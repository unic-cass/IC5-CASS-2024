* NGSPICE file created from lovers_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

.subckt lovers_controller becStatus[0] becStatus[1] becStatus[2] becStatus[3] data_in[0]
+ data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7]
+ data_in[8] data_in[9] data_out[0] data_out[10] data_out[11] data_out[12] data_out[13]
+ data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[1]
+ data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26]
+ data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] io_oeb io_out
+ ki la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7]
+ la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3]
+ la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ load_data load_status[0] load_status[1] load_status[2] load_status[3] load_status[4]
+ load_status[5] next_key slv_done slv_enable vccd1 vssd1 wb_clk_i wb_rst_i
XFILLER_0_193_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _18292_/Q _16381_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _09015_/A hold432/X vssd1 vssd1 vccd1 vccd1 _15933_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08553_ _12418_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _15900_/D sky130_fd_sc_hd__and2_1
XFILLER_0_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08484_ _14878_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ hold2630/X _09106_/B _09104_/Y _12975_/A vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09036_ hold568/X hold632/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold340 hold340/A vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 hold55/X vssd1 vssd1 vccd1 vccd1 input17/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold373 hold373/A vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold384 hold384/A vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold395 hold395/A vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _15026_/A vssd1 vssd1 vccd1 vccd1 _15204_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout831 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__buf_4
Xfanout842 _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/C1 sky130_fd_sc_hd__buf_4
X_09938_ hold3207/X hold5054/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__mux2_1
Xfanout853 _15217_/A vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__clkbuf_16
Xfanout864 fanout873/X vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__clkbuf_8
Xfanout875 _14862_/A vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__buf_8
Xfanout886 _15195_/A vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__buf_12
X_09869_ hold1466/X hold4709/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__mux2_1
Xfanout897 _14974_/A vssd1 vssd1 vccd1 vccd1 _14116_/A sky130_fd_sc_hd__buf_12
Xhold1040 _15696_/Q vssd1 vssd1 vccd1 vccd1 hold1040/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1051 _09191_/X vssd1 vssd1 vccd1 vccd1 _16207_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1062 _08453_/X vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ hold1737/X _17124_/Q _12029_/S vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__mux2_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1073 _15023_/X vssd1 vssd1 vccd1 vccd1 _15024_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_25_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_25_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ hold2221/X hold3145/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_212_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1084 hold1136/X vssd1 vssd1 vccd1 vccd1 hold1084/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _14813_/X vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11831_ hold2671/X hold4787/X _13862_/C vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14550_ hold2943/X _14535_/B _14549_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _14550_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _17078_/Q _11762_/B _11762_/C vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and3_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13501_ hold4251/X _13883_/B _13500_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13501_/X
+ sky130_fd_sc_hd__o211a_1
X_10713_ _11100_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14946_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nand2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ hold2838/X hold5595/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_344_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17749_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _17455_/CLK _16220_/D vssd1 vssd1 vccd1 vccd1 _16220_/Q sky130_fd_sc_hd__dfxtp_1
X_13432_ hold3848/X _13814_/B _13431_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10644_ hold3575/X _10998_/A _10643_/X vssd1 vssd1 vccd1 vccd1 _10644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16151_ _17508_/CLK _16151_/D vssd1 vssd1 vccd1 vccd1 _16151_/Q sky130_fd_sc_hd__dfxtp_1
X_10575_ hold4606/X _11082_/A _10574_/X vssd1 vssd1 vccd1 vccd1 _10575_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ hold4465/X _13847_/B _13362_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ hold5984/X _15113_/B hold383/X _15058_/A vssd1 vssd1 vccd1 vccd1 hold384/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12314_ _17262_/Q _12314_/B _12314_/C vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and3_1
X_16082_ _18404_/CLK _16082_/D vssd1 vssd1 vccd1 vccd1 hold832/A sky130_fd_sc_hd__dfxtp_1
X_13294_ _13294_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15033_ _14910_/A hold2507/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ hold2969/X hold4417/X _12365_/C vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ hold1523/X hold3478/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ _11694_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16984_ _17862_/CLK _16984_/D vssd1 vssd1 vccd1 vccd1 _16984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15935_ _17315_/CLK _15935_/D vssd1 vssd1 vccd1 vccd1 hold586/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11058_ _11136_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__or2_1
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18045_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10009_ _11203_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _16493_/D sky130_fd_sc_hd__nor2_1
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _17681_/CLK _15866_/D vssd1 vssd1 vccd1 vccd1 _15866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ hold1839/X _14828_/B _14816_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14817_/X
+ sky130_fd_sc_hd__o211a_1
X_17605_ _17701_/CLK _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _17696_/CLK _15797_/D vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17536_ _18364_/CLK _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14748_ _14910_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ _17479_/CLK _17467_/D vssd1 vssd1 vccd1 vccd1 _17467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14679_ hold2787/X _14666_/B _14678_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ _18391_/CLK _16418_/D vssd1 vssd1 vccd1 vccd1 _16418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ _18450_/CLK _17398_/D vssd1 vssd1 vccd1 vccd1 _17398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ _18292_/CLK _16349_/D vssd1 vssd1 vccd1 vccd1 _16349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6007 hold6035/X vssd1 vssd1 vccd1 vccd1 hold6007/X sky130_fd_sc_hd__buf_1
Xhold6018 _17523_/Q vssd1 vssd1 vccd1 vccd1 hold6018/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6029 _18409_/Q vssd1 vssd1 vccd1 vccd1 hold6029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5306 _17139_/Q vssd1 vssd1 vccd1 vccd1 hold5306/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5317 _10201_/X vssd1 vssd1 vccd1 vccd1 _16557_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5328 _17267_/Q vssd1 vssd1 vccd1 vccd1 hold5328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5339 _11464_/X vssd1 vssd1 vccd1 vccd1 _16978_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4605 _10065_/Y vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _18019_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4616 hold6046/X vssd1 vssd1 vccd1 vccd1 hold4616/X sky130_fd_sc_hd__clkbuf_2
Xhold4627 _16525_/Q vssd1 vssd1 vccd1 vccd1 hold4627/X sky130_fd_sc_hd__buf_2
XFILLER_0_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4638 _10608_/Y vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4649 _16543_/Q vssd1 vssd1 vccd1 vccd1 hold4649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3904 _16988_/Q vssd1 vssd1 vccd1 vccd1 hold3904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3915 _10999_/X vssd1 vssd1 vccd1 vccd1 _16823_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3926 _16817_/Q vssd1 vssd1 vccd1 vccd1 hold3926/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3937 _09841_/X vssd1 vssd1 vccd1 vccd1 _16437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3948 _16937_/Q vssd1 vssd1 vccd1 vccd1 hold3948/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3959 _10453_/X vssd1 vssd1 vccd1 vccd1 _16641_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout149 _12749_/S vssd1 vssd1 vccd1 vccd1 _12755_/S sky130_fd_sc_hd__buf_4
XFILLER_0_226_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07984_ _15553_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07984_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09723_ _09963_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _09960_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ hold113/X hold628/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08606_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09585_ _10560_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ hold215/X hold258/X _08536_/S vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__mux2_1
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08467_ hold5999/X _08488_/B _08466_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08398_ hold1223/X _08440_/A2 _08397_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _08398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ hold4065/X _10622_/B _10359_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _12418_/A hold724/X vssd1 vssd1 vccd1 vccd1 _16126_/D sky130_fd_sc_hd__and2_1
Xhold5840 _18398_/Q vssd1 vssd1 vccd1 vccd1 hold5840/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10291_ hold3716/X _10577_/B _10290_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10291_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5851 hold6007/X vssd1 vssd1 vccd1 vccd1 hold5851/X sky130_fd_sc_hd__clkbuf_2
Xhold5862 hold960/X vssd1 vssd1 vccd1 vccd1 hold5862/X sky130_fd_sc_hd__buf_1
XFILLER_0_143_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5873 _18416_/Q vssd1 vssd1 vccd1 vccd1 hold5873/X sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ _12261_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__or2_1
Xhold5884 hold5884/A vssd1 vssd1 vccd1 vccd1 hold5884/X sky130_fd_sc_hd__clkbuf_4
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5895 _18423_/Q vssd1 vssd1 vccd1 vccd1 hold5895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__clkbuf_8
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout650 _12804_/A vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout661 _15502_/A vssd1 vssd1 vccd1 vccd1 _15500_/A sky130_fd_sc_hd__buf_4
Xfanout672 fanout692/X vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__buf_4
Xfanout683 _14554_/C1 vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__buf_4
X_13981_ hold2319/X _13986_/B _13980_/Y _13921_/A vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout694 _12600_/A vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__buf_4
XFILLER_0_38_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15720_ _17221_/CLK _15720_/D vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ hold3251/X _12931_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__mux2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _17195_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ hold3297/X _12862_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14602_ _15103_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__or2_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18370_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11814_ _12288_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15582_ _17639_/CLK _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ hold3177/X _12793_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12794_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_205_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17321_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _17321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _15105_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__or2_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ hold3567/X _11652_/A _11744_/X vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17252_ _17897_/CLK _17252_/D vssd1 vssd1 vccd1 vccd1 _17252_/Q sky130_fd_sc_hd__dfxtp_1
X_14464_ hold1682/X _14482_/A2 _14463_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14464_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11676_ _12243_/A _11676_/B vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__or2_1
X_16203_ _17435_/CLK _16203_/D vssd1 vssd1 vccd1 vccd1 _16203_/Q sky130_fd_sc_hd__dfxtp_1
X_13415_ hold1223/X _17592_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13416_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10627_ _18461_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _16699_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17183_ _17215_/CLK _17183_/D vssd1 vssd1 vccd1 vccd1 _17183_/Q sky130_fd_sc_hd__dfxtp_1
X_14395_ _14968_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _17329_/CLK _16134_/D vssd1 vssd1 vccd1 vccd1 hold616/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ hold2029/X hold5663/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10558_ hold3695/X _11192_/B _10557_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _16676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ _18410_/CLK _16065_/D vssd1 vssd1 vccd1 vccd1 hold396/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13277_ _13276_/X hold4649/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10489_ hold4980/X _10601_/B _10488_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ hold719/X _15016_/B vssd1 vssd1 vccd1 vccd1 hold720/A sky130_fd_sc_hd__or2_1
XFILLER_0_227_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12228_ _12234_/A _12228_/B vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _12231_/A _12159_/B vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1809 _17833_/Q vssd1 vssd1 vccd1 vccd1 hold1809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16967_ _18427_/CLK _16967_/D vssd1 vssd1 vccd1 vccd1 _16967_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _16081_/CLK _15918_/D vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16898_ _17971_/CLK _16898_/D vssd1 vssd1 vccd1 vccd1 _16898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ _17734_/CLK _15849_/D vssd1 vssd1 vccd1 vccd1 _15849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_266_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18055_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09370_ hold586/X _15486_/A2 _15488_/A2 hold584/X vssd1 vssd1 vccd1 vccd1 _09370_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ _15545_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17519_ _17525_/CLK _17519_/D vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08252_ _14758_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _14403_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5103 _11760_/Y vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5114 _17169_/Q vssd1 vssd1 vccd1 vccd1 hold5114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5125 _11494_/X vssd1 vssd1 vccd1 vccd1 _16988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5136 _16638_/Q vssd1 vssd1 vccd1 vccd1 hold5136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4402 _11989_/X vssd1 vssd1 vccd1 vccd1 _17153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5147 _11908_/X vssd1 vssd1 vccd1 vccd1 _17126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4413 _17643_/Q vssd1 vssd1 vccd1 vccd1 hold4413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5158 _17069_/Q vssd1 vssd1 vccd1 vccd1 hold5158/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5169 _10801_/X vssd1 vssd1 vccd1 vccd1 _16757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4424 _12175_/X vssd1 vssd1 vccd1 vccd1 _17215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4435 _17207_/Q vssd1 vssd1 vccd1 vccd1 hold4435/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3701 _17394_/Q vssd1 vssd1 vccd1 vccd1 hold3701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4446 _11893_/X vssd1 vssd1 vccd1 vccd1 _17121_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3712 _16563_/Q vssd1 vssd1 vccd1 vccd1 hold3712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4457 _16839_/Q vssd1 vssd1 vccd1 vccd1 hold4457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3723 _11775_/Y vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4468 _11017_/X vssd1 vssd1 vccd1 vccd1 _16829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4479 _17739_/Q vssd1 vssd1 vccd1 vccd1 hold4479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3734 _17119_/Q vssd1 vssd1 vccd1 vccd1 hold3734/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3745 _10228_/X vssd1 vssd1 vccd1 vccd1 _16566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3756 _17404_/Q vssd1 vssd1 vccd1 vccd1 hold3756/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3767 _10528_/X vssd1 vssd1 vccd1 vccd1 _16666_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3778 _17434_/Q vssd1 vssd1 vccd1 vccd1 hold3778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3789 _16570_/Q vssd1 vssd1 vccd1 vccd1 hold3789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07967_ hold1294/X _07978_/B _07966_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _07967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ hold4059/X _10013_/B _09705_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07898_ _15521_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07898_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09637_ hold4000/X _10010_/B _09636_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09637_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09568_ hold4735/X _10049_/B _09567_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09568_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08519_ _17523_/Q _17522_/Q vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09499_ _18459_/Q _12510_/B vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ hold5216/X _11617_/A2 _11529_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11530_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ hold4493/X _12314_/B _11460_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13193_/X _13199_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17543_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_163_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10412_ hold1344/X _16628_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ hold5505/X _12338_/B _11391_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11392_/X
+ sky130_fd_sc_hd__o211a_1
X_14180_ _15199_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13130_/X hold4674/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__mux2_1
X_10343_ hold2260/X hold4970/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5670 _09580_/X vssd1 vssd1 vccd1 vccd1 _16350_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10274_ hold1964/X hold4131/X _10580_/C vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__mux2_1
X_13062_ _13062_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__or2_1
Xhold5681 _17568_/Q vssd1 vssd1 vccd1 vccd1 hold5681/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5692 _13672_/X vssd1 vssd1 vccd1 vccd1 _17677_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12013_ hold5156/X _12299_/B _12012_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _12013_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4980 _16685_/Q vssd1 vssd1 vccd1 vccd1 hold4980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17870_ _17870_/CLK _17870_/D vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4991 _11431_/X vssd1 vssd1 vccd1 vccd1 _16967_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16821_ _18054_/CLK _16821_/D vssd1 vssd1 vccd1 vccd1 _16821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout480 _11219_/C vssd1 vssd1 vccd1 vccd1 _11789_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout491 _10019_/C vssd1 vssd1 vccd1 vccd1 _10010_/C sky130_fd_sc_hd__buf_6
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16752_ _17985_/CLK _16752_/D vssd1 vssd1 vccd1 vccd1 _16752_/Q sky130_fd_sc_hd__dfxtp_1
X_13964_ _15525_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _17775_/CLK _15703_/D vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfxtp_1
X_12915_ _12921_/A _12915_/B vssd1 vssd1 vccd1 vccd1 _17481_/D sky130_fd_sc_hd__and2_1
X_16683_ _18294_/CLK _16683_/D vssd1 vssd1 vccd1 vccd1 _16683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _15496_/A _13895_/B vssd1 vssd1 vccd1 vccd1 _17753_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18422_ _18422_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _17166_/CLK _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _12870_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _17458_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18353_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _17900_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12780_/A _12777_/B vssd1 vssd1 vccd1 vccd1 _17435_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17304_ _17304_/CLK _17304_/D vssd1 vssd1 vccd1 vccd1 hold788/A sky130_fd_sc_hd__dfxtp_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14516_ hold2577/X _14535_/B _14515_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14516_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _18356_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11728_ _12310_/A _11728_/B vssd1 vssd1 vccd1 vccd1 _17066_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_232_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15496_ _15496_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17235_ _17899_/CLK _17235_/D vssd1 vssd1 vccd1 vccd1 _17235_/Q sky130_fd_sc_hd__dfxtp_1
X_14447_ _15128_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_226_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11659_ hold5577/X _11753_/B _11658_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ _17166_/CLK _17166_/D vssd1 vssd1 vccd1 vccd1 _17166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14378_ _14378_/A hold427/X vssd1 vssd1 vccd1 vccd1 _17986_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold906 hold906/A vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold917 becStatus[2] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ _17340_/CLK _16117_/D vssd1 vssd1 vccd1 vccd1 _16117_/Q sky130_fd_sc_hd__dfxtp_1
Xhold928 hold928/A vssd1 vssd1 vccd1 vccd1 hold928/X sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _13713_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__or2_1
Xhold939 hold939/A vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _17129_/CLK _17097_/D vssd1 vssd1 vccd1 vccd1 _17097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _17304_/CLK _16048_/D vssd1 vssd1 vccd1 vccd1 hold652/A sky130_fd_sc_hd__dfxtp_1
Xhold3008 _18377_/Q vssd1 vssd1 vccd1 vccd1 hold3008/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3019 _15836_/Q vssd1 vssd1 vccd1 vccd1 hold3019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2307 _14015_/X vssd1 vssd1 vccd1 vccd1 _17811_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08870_ hold554/X hold661/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__mux2_1
XFILLER_0_110_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2318 _14247_/X vssd1 vssd1 vccd1 vccd1 _17922_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2329 _17889_/Q vssd1 vssd1 vccd1 vccd1 hold2329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07821_ _15555_/A _15551_/A _15553_/A vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__or3b_1
Xhold1606 _08257_/X vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1617 _14191_/X vssd1 vssd1 vccd1 vccd1 _17896_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1628 _15737_/Q vssd1 vssd1 vccd1 vccd1 hold1628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17999_ _17999_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1639 _14973_/X vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_447_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17623_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_224_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09422_ _09438_/B _16297_/Q vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09353_ _15547_/A hold181/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__or3_2
XFILLER_0_158_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08304_ hold2373/X _08336_/A2 _08303_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09284_ _12780_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _16253_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08235_ hold1674/X _08263_/A2 _08234_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08166_ _15517_/A hold2019/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08097_ hold2384/X _08097_/A2 _08096_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _08097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4210 _13708_/X vssd1 vssd1 vccd1 vccd1 _17689_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4221 _17149_/Q vssd1 vssd1 vccd1 vccd1 hold4221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4232 _15293_/X vssd1 vssd1 vccd1 vccd1 _15294_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4243 _17641_/Q vssd1 vssd1 vccd1 vccd1 hold4243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4254 _11998_/X vssd1 vssd1 vccd1 vccd1 _17156_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3520 _13600_/X vssd1 vssd1 vccd1 vccd1 _17653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4265 _17068_/Q vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3531 _17672_/Q vssd1 vssd1 vccd1 vccd1 hold3531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4276 _11446_/X vssd1 vssd1 vccd1 vccd1 _16972_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3542 _09388_/X vssd1 vssd1 vccd1 vccd1 _16282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4287 _17734_/Q vssd1 vssd1 vccd1 vccd1 hold4287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3553 _16527_/Q vssd1 vssd1 vccd1 vccd1 hold3553/X sky130_fd_sc_hd__buf_2
Xhold4298 _13489_/X vssd1 vssd1 vccd1 vccd1 _17616_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3564 _11727_/Y vssd1 vssd1 vccd1 vccd1 _11728_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2830 _18101_/Q vssd1 vssd1 vccd1 vccd1 hold2830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3575 _16545_/Q vssd1 vssd1 vccd1 vccd1 hold3575/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3586 _17360_/Q vssd1 vssd1 vccd1 vccd1 hold3586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 _14540_/X vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 _18173_/Q vssd1 vssd1 vccd1 vccd1 hold2852/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _13046_/C _12445_/B vssd1 vssd1 vccd1 vccd1 _09006_/S sky130_fd_sc_hd__or2_2
XFILLER_0_214_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3597 _12348_/Y vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2863 _14801_/X vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_188_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18360_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2874 _18017_/Q vssd1 vssd1 vccd1 vccd1 hold2874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 _14599_/X vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2896 _15790_/Q vssd1 vssd1 vccd1 vccd1 hold2896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_117_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17313_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ hold911/X hold5471/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ hold2765/X hold3779/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13680_ _13776_/A _13680_/B vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ hold1129/X hold4753/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ hold2136/X hold3336/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15350_ hold907/X _09367_/A _09392_/A hold891/X vssd1 vssd1 vccd1 vccd1 _15350_/X
+ sky130_fd_sc_hd__a22o_1
X_12562_ hold1090/X hold3472/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ hold2957/X hold756/X _14300_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14301_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11513_ _17841_/Q hold4439/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__mux2_1
X_15281_ _16292_/Q _15477_/A2 _15487_/B1 hold156/X _15280_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/D sky130_fd_sc_hd__a221o_1
X_12493_ hold62/X _12509_/A2 _12507_/A3 _12492_/X _12444_/A vssd1 vssd1 vccd1 vccd1
+ hold63/A sky130_fd_sc_hd__o311a_1
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17020_ _17898_/CLK _17020_/D vssd1 vssd1 vccd1 vccd1 _17020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14232_ _14913_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__nor2_1
X_11444_ hold1656/X _16972_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14843_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14206_/B sky130_fd_sc_hd__or2_4
XFILLER_0_225_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ hold2319/X _16949_/Q _11768_/C vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _17565_/Q _17099_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_237_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10326_ _10542_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__or2_1
X_14094_ _15547_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__nand2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _17524_/Q hold933/X _13044_/X _13056_/C _13048_/A vssd1 vssd1 vccd1 vccd1
+ hold934/A sky130_fd_sc_hd__o221a_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _17952_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_1
X_10257_ _10998_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10257_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10188_ _10533_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__or2_1
X_17853_ _17885_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16804_ _18071_/CLK _16804_/D vssd1 vssd1 vccd1 vccd1 _16804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14996_ _15103_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__or2_1
X_17784_ _17816_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16735_ _17960_/CLK _16735_/D vssd1 vssd1 vccd1 vccd1 _16735_/Q sky130_fd_sc_hd__dfxtp_1
X_13947_ _14627_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _13996_/B sky130_fd_sc_hd__or2_4
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _18222_/CLK _16666_/D vssd1 vssd1 vccd1 vccd1 _16666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ hold3740/X _13782_/A _13877_/X vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18405_ _18405_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15617_ _17273_/CLK _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ hold2186/X _17454_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__mux2_1
X_16597_ _18199_/CLK _16597_/D vssd1 vssd1 vccd1 vccd1 _16597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18336_ _18366_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
X_15548_ hold2361/X _15547_/B _15547_/Y _15548_/C1 vssd1 vssd1 vccd1 vccd1 _15548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18267_ _18375_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _17323_/Q _09357_/A _15479_/B1 _16024_/Q _15478_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08020_ hold2719/X _08029_/B _08019_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _08020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17218_ _17639_/CLK _17218_/D vssd1 vssd1 vccd1 vccd1 _17218_/Q sky130_fd_sc_hd__dfxtp_1
X_18198_ _18198_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold714 hold714/A vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17149_ _17273_/CLK _17149_/D vssd1 vssd1 vccd1 vccd1 _17149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 hold725/A vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/A vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 hold758/A vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09971_ _18392_/Q hold3681/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__mux2_1
Xhold769 hold769/A vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ hold210/X hold464/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold465/A sky130_fd_sc_hd__mux2_1
Xhold2104 _17799_/Q vssd1 vssd1 vccd1 vccd1 hold2104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _18200_/Q vssd1 vssd1 vccd1 vccd1 hold2115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 _12974_/X vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ _12416_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _16045_/D sky130_fd_sc_hd__and2_1
Xhold2137 _15522_/X vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _14512_/X vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _14077_/X vssd1 vssd1 vccd1 vccd1 _17841_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _08418_/X vssd1 vssd1 vccd1 vccd1 _15839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _15745_/Q vssd1 vssd1 vccd1 vccd1 hold1414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1425 _15611_/Q vssd1 vssd1 vccd1 vccd1 hold1425/X sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ _07804_/A _16286_/Q vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__and2_2
XFILLER_0_139_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_281_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18200_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1436 _15585_/Q vssd1 vssd1 vccd1 vccd1 hold1436/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1447 _14113_/X vssd1 vssd1 vccd1 vccd1 _17858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08784_ _15482_/A hold211/X vssd1 vssd1 vccd1 vccd1 _16012_/D sky130_fd_sc_hd__and2_1
Xhold1458 _17963_/Q vssd1 vssd1 vccd1 vccd1 hold1458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _14179_/X vssd1 vssd1 vccd1 vccd1 _17890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_210_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ _07804_/A hold5916/X _15264_/A _09404_/X vssd1 vssd1 vccd1 vccd1 _09405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ hold1877/X _09338_/A2 _09335_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09267_ hold246/A _16245_/Q _09273_/S vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08218_ hold1414/X _08213_/B _08217_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08218_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ hold944/X _09220_/B vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ _08149_/A _08149_/B vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__and2_1
XFILLER_0_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ hold4666/X _11064_/A _11159_/X vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4040 _16497_/Q vssd1 vssd1 vccd1 vccd1 hold4040/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10111_ hold4936/X _10477_/A2 _10110_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10111_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4051 _09910_/X vssd1 vssd1 vccd1 vccd1 _16460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4062 _10411_/X vssd1 vssd1 vccd1 vccd1 _16627_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _11103_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11091_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_369_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4073 _17660_/Q vssd1 vssd1 vccd1 vccd1 hold4073/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4084 _13513_/X vssd1 vssd1 vccd1 vccd1 _17624_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3350 _09805_/X vssd1 vssd1 vccd1 vccd1 _16425_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4095 _16853_/Q vssd1 vssd1 vccd1 vccd1 hold4095/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3361 _16361_/Q vssd1 vssd1 vccd1 vccd1 hold3361/X sky130_fd_sc_hd__dlygate4sd3_1
X_10042_ _11194_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _16504_/D sky130_fd_sc_hd__nor2_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3372 _17417_/Q vssd1 vssd1 vccd1 vccd1 hold3372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3383 _17481_/Q vssd1 vssd1 vccd1 vccd1 hold3383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__buf_4
XFILLER_0_227_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3394 _17476_/Q vssd1 vssd1 vccd1 vccd1 hold3394/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2660 _15779_/Q vssd1 vssd1 vccd1 vccd1 hold2660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _15189_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__or2_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2671 _15693_/Q vssd1 vssd1 vccd1 vccd1 hold2671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__buf_4
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2682 _14408_/X vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2693 _18068_/Q vssd1 vssd1 vccd1 vccd1 hold2693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ hold4114/X _13814_/B _13800_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _17720_/D
+ sky130_fd_sc_hd__o211a_1
Xhold1970 _18227_/Q vssd1 vssd1 vccd1 vccd1 hold1970/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1981 _18260_/Q vssd1 vssd1 vccd1 vccd1 hold1981/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ hold2915/X _14772_/B _14780_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14781_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1992 _15732_/Q vssd1 vssd1 vccd1 vccd1 hold1992/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ hold2192/X hold4342/X _13877_/C vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__mux2_1
X_16520_ _18112_/CLK _16520_/D vssd1 vssd1 vccd1 vccd1 _16520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13732_ hold5715/X _13832_/B _13731_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13732_/X
+ sky130_fd_sc_hd__o211a_1
X_10944_ _11136_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16451_ _18266_/CLK _16451_/D vssd1 vssd1 vccd1 vccd1 _16451_/Q sky130_fd_sc_hd__dfxtp_1
X_13663_ hold4185/X _13883_/B _13662_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13663_/X
+ sky130_fd_sc_hd__o211a_1
X_10875_ _11106_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__or2_1
X_15402_ _15480_/A _15402_/B _15402_/C _15402_/D vssd1 vssd1 vccd1 vccd1 _15402_/X
+ sky130_fd_sc_hd__or4_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12614_ hold3292/X _12613_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _18293_/CLK _16382_/D vssd1 vssd1 vccd1 vccd1 _16382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13594_ hold4372/X _13880_/B _13593_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13594_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18193_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15333_ _15490_/A1 _15325_/X _15332_/X _15490_/B1 _18407_/Q vssd1 vssd1 vccd1 vccd1
+ _15333_/X sky130_fd_sc_hd__a32o_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12545_ hold3557/X _12544_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17257_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _18052_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ _15264_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__and2_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12476_ _17331_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ _17975_/CLK _17003_/D vssd1 vssd1 vccd1 vccd1 _17003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14215_ hold1825/X _14198_/B _14214_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14215_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_5 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _11712_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
X_15195_ _15195_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14146_ _15545_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nand2_1
X_11358_ _12219_/A _11358_/B vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10309_ hold4938/X _10619_/B _10308_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14077_ hold6008/X _14107_/A2 _14076_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11289_ _11694_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _13029_/B hold958/X _13028_/C vssd1 vssd1 vccd1 vccd1 _17519_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_225_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17905_ _17905_/CLK _17905_/D vssd1 vssd1 vccd1 vccd1 _17905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _17867_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _17767_/CLK _17767_/D vssd1 vssd1 vccd1 vccd1 _17767_/Q sky130_fd_sc_hd__dfxtp_1
X_14979_ hold5998/X hold514/X _14978_/X _15044_/A vssd1 vssd1 vccd1 vccd1 hold515/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16718_ _18060_/CLK _16718_/D vssd1 vssd1 vccd1 vccd1 _16718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17698_ _17730_/CLK _17698_/D vssd1 vssd1 vccd1 vccd1 _17698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16649_ _18201_/CLK _16649_/D vssd1 vssd1 vccd1 vccd1 _16649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _15555_/A _09121_/B _15553_/A _15551_/A vssd1 vssd1 vccd1 vccd1 _09400_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18319_ _18319_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09052_ hold210/X hold232/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08003_ _14403_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold500 hold556/X vssd1 vssd1 vccd1 vccd1 hold557/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold511 hold751/X vssd1 vssd1 vccd1 vccd1 hold752/A sky130_fd_sc_hd__buf_4
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold533 hold533/A vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__buf_6
Xhold544 hold544/A vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold555 hold555/A vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 hold82/X vssd1 vssd1 vccd1 vccd1 input14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 input21/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__buf_1
Xhold588 hold588/A vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_462_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08905_ _12416_/A hold380/X vssd1 vssd1 vccd1 vccd1 _16070_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _11064_/A _09885_/B vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__or2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _08010_/X vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _14013_/X vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ hold256/X hold387/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08837_/B sky130_fd_sc_hd__mux2_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _07943_/X vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _15122_/X vssd1 vssd1 vccd1 vccd1 _18343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 _08051_/X vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1255 _09413_/X vssd1 vssd1 vccd1 vccd1 _16292_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_15_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_15_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 _13991_/X vssd1 vssd1 vccd1 vccd1 _17800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08767_ hold568/X _16004_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold569/A sky130_fd_sc_hd__mux2_1
Xhold1277 input40/X vssd1 vssd1 vccd1 vccd1 hold1277/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _13997_/X vssd1 vssd1 vccd1 vccd1 _17803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _14857_/X vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _12436_/A _08698_/B vssd1 vssd1 vccd1 vccd1 _15970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10660_ hold4211/X _11729_/B _10659_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _10660_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _15541_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ _18461_/A _10591_/B vssd1 vssd1 vccd1 vccd1 _16687_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ hold4695/X _12234_/A _12329_/X vssd1 vssd1 vccd1 vccd1 _12330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ _14681_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__nor2_1
X_11212_ _12340_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _16894_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_121_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12192_ _13716_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__or2_1
Xclkbuf_6_54_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_54_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11143_ _11158_/A _11143_/B vssd1 vssd1 vccd1 vccd1 _16871_/D sky130_fd_sc_hd__nor2_1
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 _13153_/A vssd1 vssd1 vccd1 vccd1 output75/X sky130_fd_sc_hd__buf_6
Xoutput86 _13233_/A vssd1 vssd1 vccd1 vccd1 output86/X sky130_fd_sc_hd__buf_6
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_132_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16097_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput97 _13081_/A vssd1 vssd1 vccd1 vccd1 output97/X sky130_fd_sc_hd__buf_6
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15951_ _17298_/CLK _15951_/D vssd1 vssd1 vccd1 vccd1 hold872/A sky130_fd_sc_hd__dfxtp_1
X_11074_ hold5403/X _11732_/B _11073_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _11074_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3180 _12827_/X vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10025_ _16499_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__and3_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3191 _18277_/Q vssd1 vssd1 vccd1 vccd1 hold3191/X sky130_fd_sc_hd__dlygate4sd3_1
X_14902_ _14972_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__or2_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _17254_/CLK _15882_/D vssd1 vssd1 vccd1 vccd1 _15882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2490 _18258_/Q vssd1 vssd1 vccd1 vccd1 hold2490/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _17650_/CLK _17621_/D vssd1 vssd1 vccd1 vccd1 _17621_/Q sky130_fd_sc_hd__dfxtp_1
X_14833_ hold1831/X _14828_/B _14832_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14833_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _18221_/CLK _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
X_14764_ _15103_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14764_/X sky130_fd_sc_hd__or2_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _12231_/A _11976_/B vssd1 vssd1 vccd1 vccd1 _11976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _18390_/CLK _16503_/D vssd1 vssd1 vccd1 vccd1 _16503_/Q sky130_fd_sc_hd__dfxtp_1
X_13715_ hold2564/X hold4988/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ hold5447/X _11198_/B _10926_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10927_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17483_ _17483_/CLK _17483_/D vssd1 vssd1 vccd1 vccd1 _17483_/Q sky130_fd_sc_hd__dfxtp_1
X_14695_ hold2689/X _14714_/B _14694_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16434_ _18377_/CLK _16434_/D vssd1 vssd1 vccd1 vccd1 _16434_/Q sky130_fd_sc_hd__dfxtp_1
X_13646_ hold1190/X _17669_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13647_/B sky130_fd_sc_hd__mux2_1
X_10858_ hold4387/X _11147_/B _10857_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10858_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _18276_/CLK _16365_/D vssd1 vssd1 vccd1 vccd1 _16365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ hold2660/X _17646_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13578_/B sky130_fd_sc_hd__mux2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10789_ hold4018/X _11168_/B _10788_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ _17335_/Q _15448_/B1 _15485_/B1 hold196/X vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__a22o_1
X_18104_ _18234_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ _12531_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _17352_/D sky130_fd_sc_hd__and2_1
X_16296_ _16323_/CLK _16296_/D vssd1 vssd1 vccd1 vccd1 _16296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15247_ hold288/X _15487_/A2 _15484_/B1 hold620/X _15246_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/B sky130_fd_sc_hd__a221o_1
X_18035_ _18035_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12459_ hold47/X _12509_/A2 _12507_/A3 _12458_/X _09053_/A vssd1 vssd1 vccd1 vccd1
+ hold48/A sky130_fd_sc_hd__o311a_1
Xhold4809 _16372_/Q vssd1 vssd1 vccd1 vccd1 hold4809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15178_ hold1835/X _15165_/B _15177_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15178_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ hold2345/X _14148_/B _14128_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14129_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout309 _11097_/A vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__buf_4
XFILLER_0_158_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ hold5675/X _10070_/B _09669_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08621_ hold361/X hold431/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold432/A sky130_fd_sc_hd__mux2_1
XFILLER_0_234_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17819_ _17851_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08552_ hold98/X hold867/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08483_ hold2325/X _08488_/B _08482_/Y _08137_/A vssd1 vssd1 vccd1 vccd1 _08483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09104_ _15545_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09035_ _12436_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _16134_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 hold341/A vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 input17/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__buf_1
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 hold374/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold385 hold385/A vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold396 hold396/A vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _15192_/C1 vssd1 vssd1 vccd1 vccd1 _15198_/C1 sky130_fd_sc_hd__buf_4
Xfanout821 fanout847/X vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__buf_4
X_09937_ _10031_/A _10007_/B _09936_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09937_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout832 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__buf_4
Xfanout843 fanout847/X vssd1 vssd1 vccd1 vccd1 _14849_/C1 sky130_fd_sc_hd__buf_4
Xfanout854 _07782_/Y vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__buf_8
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout865 fanout873/X vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__buf_8
Xfanout876 hold944/X vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__clkbuf_16
X_09868_ hold5090/X _10034_/B _09867_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09868_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout887 hold1029/X vssd1 vssd1 vccd1 vccd1 hold1030/A sky130_fd_sc_hd__buf_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 hold1030/A vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__buf_12
Xfanout898 hold1334/X vssd1 vssd1 vccd1 vccd1 hold1335/A sky130_fd_sc_hd__buf_6
Xhold1041 _08114_/X vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _12531_/A hold787/X vssd1 vssd1 vccd1 vccd1 _16028_/D sky130_fd_sc_hd__and2_1
Xhold1052 _16203_/Q vssd1 vssd1 vccd1 vccd1 hold1052/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _16154_/Q vssd1 vssd1 vccd1 vccd1 hold1063/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 _18326_/Q vssd1 vssd1 vccd1 vccd1 hold1074/X sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ hold3768/X _10010_/B _09798_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09799_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 hold1085/A vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__buf_12
XFILLER_0_77_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1096 _15751_/Q vssd1 vssd1 vccd1 vccd1 hold1096/X sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ hold5024/X _12308_/B _11829_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _12367_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _17077_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13788_/A _13500_/B vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__or2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ hold1636/X hold4625/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__mux2_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14480_ hold2919/X _14482_/A2 _14479_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ hold5531/X _12329_/B _11691_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11692_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13431_ _13623_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__or2_1
X_10643_ _16705_/Q _10646_/B _10997_/S vssd1 vssd1 vccd1 vccd1 _10643_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _17508_/CLK _16150_/D vssd1 vssd1 vccd1 vccd1 _16150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13362_ _13746_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10574_ _16682_/Q _11192_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__and3_1
XFILLER_0_90_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15101_ hold382/X _15125_/B vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__or2_1
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12313_ _13825_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _17261_/D sky130_fd_sc_hd__nor2_1
X_16081_ _16081_/CLK _16081_/D vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_384_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17166_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _13292_/X hold3575/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_84_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15032_ _15032_/A _15032_/B vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__and2_1
X_12244_ hold5511/X _12338_/B _12243_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _12244_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_313_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ hold4423/X _12274_/A2 _12174_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ hold1532/X _16866_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16983_ _17902_/CLK _16983_/D vssd1 vssd1 vccd1 vccd1 _16983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15934_ _18411_/CLK _15934_/D vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__dfxtp_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ hold1968/X _16843_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10008_ _13134_/A _09936_/A _10007_/X vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _17738_/CLK _15865_/D vssd1 vssd1 vccd1 vccd1 _15865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _17680_/CLK _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
X_14816_ _15209_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _17730_/CLK _15796_/D vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _18364_/CLK _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14747_ hold2812/X _14774_/B _14746_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ hold4485/X _12365_/B _11958_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _15233_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14678_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _17479_/CLK _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16417_ _16517_/CLK _16417_/D vssd1 vssd1 vccd1 vccd1 _16417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13629_ _13734_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__or2_1
XFILLER_0_229_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17397_ _18448_/CLK _17397_/D vssd1 vssd1 vccd1 vccd1 _17397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16348_ _18387_/CLK _16348_/D vssd1 vssd1 vccd1 vccd1 _16348_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6008 _17841_/Q vssd1 vssd1 vccd1 vccd1 hold6008/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6019 _18420_/Q vssd1 vssd1 vccd1 vccd1 hold6019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16279_ _17379_/CLK _16279_/D vssd1 vssd1 vccd1 vccd1 _16279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5307 _11851_/X vssd1 vssd1 vccd1 vccd1 _17107_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5318 _16858_/Q vssd1 vssd1 vccd1 vccd1 hold5318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5329 _12235_/X vssd1 vssd1 vccd1 vccd1 _17235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4606 _16522_/Q vssd1 vssd1 vccd1 vccd1 hold4606/X sky130_fd_sc_hd__buf_2
X_18018_ _18018_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4617 _16547_/Q vssd1 vssd1 vccd1 vccd1 hold4617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4628 _10584_/Y vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4639 _16541_/Q vssd1 vssd1 vccd1 vccd1 hold4639/X sky130_fd_sc_hd__buf_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3905 _11398_/X vssd1 vssd1 vccd1 vccd1 _16956_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3916 _16674_/Q vssd1 vssd1 vccd1 vccd1 hold3916/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3927 _10885_/X vssd1 vssd1 vccd1 vccd1 _16785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3938 _17655_/Q vssd1 vssd1 vccd1 vccd1 hold3938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3949 _11245_/X vssd1 vssd1 vccd1 vccd1 _16905_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07983_ hold1371/X _07991_/A2 _07982_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09722_ hold2676/X _16398_/Q _10034_/C vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09653_ hold1966/X hold3619/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08604_ _12412_/A hold760/X vssd1 vssd1 vccd1 vccd1 _15924_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ hold1430/X _13286_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _09055_/A hold507/X vssd1 vssd1 vccd1 vccd1 _15891_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _15199_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08397_ hold999/X _08445_/B vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5830 output83/X vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_12
X_09018_ hold163/X hold723/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold724/A sky130_fd_sc_hd__mux2_1
XFILLER_0_104_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10290_ _10482_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5841 _18401_/Q vssd1 vssd1 vccd1 vccd1 hold5841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5852 hold5852/A vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_12
Xhold5863 _16281_/Q vssd1 vssd1 vccd1 vccd1 hold5863/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5874 hold5874/A vssd1 vssd1 vccd1 vccd1 hold5874/X sky130_fd_sc_hd__clkbuf_4
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5885 hold6019/X vssd1 vssd1 vccd1 vccd1 hold5885/X sky130_fd_sc_hd__clkbuf_4
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5896 hold5896/A vssd1 vssd1 vccd1 vccd1 hold5896/X sky130_fd_sc_hd__buf_4
XFILLER_0_218_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout640 _12807_/A vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__buf_2
Xfanout651 fanout693/X vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__buf_4
Xfanout662 fanout693/X vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13980_ _14946_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_205_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout673 _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__buf_4
Xfanout684 _14554_/C1 vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__buf_4
Xfanout695 _12600_/A vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__buf_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ hold1176/X _17488_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12931_/X sky130_fd_sc_hd__mux2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15650_ _17161_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ hold1057/X _17465_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14601_ hold1797/X _14612_/B _14600_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14601_/X
+ sky130_fd_sc_hd__o211a_1
X_11813_ hold2526/X _17095_/Q _12302_/C vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__mux2_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _17217_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ hold3049/X _17442_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__mux2_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17320_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 _17320_/Q sky130_fd_sc_hd__dfxtp_1
X_14532_ hold3104/X _14535_/B _14531_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _14532_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11744_ _17072_/Q _12317_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__and3_1
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14517_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14463_/X sky130_fd_sc_hd__or2_1
X_17251_ _17283_/CLK _17251_/D vssd1 vssd1 vccd1 vccd1 _17251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11675_ hold1448/X hold4350/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13414_ hold5172/X _13798_/A2 _13413_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _13414_/X
+ sky130_fd_sc_hd__o211a_1
X_16202_ _18453_/CLK _16202_/D vssd1 vssd1 vccd1 vccd1 _16202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ hold4621/X _10533_/A _10625_/X vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17182_ _17234_/CLK _17182_/D vssd1 vssd1 vccd1 vccd1 _17182_/Q sky130_fd_sc_hd__dfxtp_1
X_14394_ hold733/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__or2_4
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _17340_/CLK _16133_/D vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13345_ hold5743/X _13832_/B _13344_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13345_/X
+ sky130_fd_sc_hd__o211a_1
X_10557_ _11100_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ _18405_/CLK _16064_/D vssd1 vssd1 vccd1 vccd1 hold891/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ hold4693/X _13275_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_122_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10488_ _10488_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10488_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15015_ hold1318/X hold514/X _15014_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15015_/X
+ sky130_fd_sc_hd__o211a_1
X_12227_ hold2182/X hold4305/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ hold1427/X _17210_/Q _13868_/C vssd1 vssd1 vccd1 vccd1 _12159_/B sky130_fd_sc_hd__mux2_1
X_11109_ _11658_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__or2_1
X_12089_ hold2905/X _17187_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16966_ _17876_/CLK _16966_/D vssd1 vssd1 vccd1 vccd1 _16966_/Q sky130_fd_sc_hd__dfxtp_1
X_15917_ _18407_/CLK _15917_/D vssd1 vssd1 vccd1 vccd1 hold158/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16897_ _17970_/CLK _16897_/D vssd1 vssd1 vccd1 vccd1 _16897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _17734_/CLK _15848_/D vssd1 vssd1 vccd1 vccd1 _15848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15779_ _17731_/CLK _15779_/D vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08320_ hold2004/X _08323_/B _08319_/Y _12657_/A vssd1 vssd1 vccd1 vccd1 _08320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _17525_/CLK _17518_/D vssd1 vssd1 vccd1 vccd1 _17518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ hold5975/X _08263_/A2 hold1303/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17449_ _17878_/CLK _17449_/D vssd1 vssd1 vccd1 vccd1 _17449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_235_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18159_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08182_ hold2557/X _08209_/B _08181_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5104 _16430_/Q vssd1 vssd1 vccd1 vccd1 hold5104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5115 _11941_/X vssd1 vssd1 vccd1 vccd1 _17137_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5126 _16680_/Q vssd1 vssd1 vccd1 vccd1 hold5126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5137 _10348_/X vssd1 vssd1 vccd1 vccd1 _16606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5148 _16762_/Q vssd1 vssd1 vccd1 vccd1 hold5148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4403 _16761_/Q vssd1 vssd1 vccd1 vccd1 hold4403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4414 _13474_/X vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5159 _11641_/X vssd1 vssd1 vccd1 vccd1 _17037_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4425 _16829_/Q vssd1 vssd1 vccd1 vccd1 hold4425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4436 _12055_/X vssd1 vssd1 vccd1 vccd1 _17175_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4447 _16012_/Q vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3702 _17574_/Q vssd1 vssd1 vccd1 vccd1 hold3702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3713 _10123_/X vssd1 vssd1 vccd1 vccd1 _16531_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4458 _10951_/X vssd1 vssd1 vccd1 vccd1 _16807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3724 _17111_/Q vssd1 vssd1 vccd1 vccd1 hold3724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4469 _17054_/Q vssd1 vssd1 vccd1 vccd1 hold4469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3735 _12366_/Y vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3746 _17029_/Q vssd1 vssd1 vccd1 vccd1 hold3746/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3757 _12683_/X vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3768 _16455_/Q vssd1 vssd1 vccd1 vccd1 hold3768/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3779 _17411_/Q vssd1 vssd1 vccd1 vccd1 hold3779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _15535_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09705_ _09918_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07897_ hold1456/X _07918_/B _07896_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _07897_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ _09933_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09567_ _09954_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08518_ hold2083/X _08503_/Y _08517_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _08518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09498_ _14681_/A _09498_/B _09498_/C _09498_/D vssd1 vssd1 vccd1 vccd1 _12510_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ hold203/X _14913_/A vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__or2_4
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _12243_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ hold4061/X _10637_/B _10410_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11391_ _12243_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ _17567_/Q _17101_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10342_ hold3954/X _10628_/B _10341_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10342_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ _13060_/X hold3695/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
Xhold5660 _13821_/Y vssd1 vssd1 vccd1 vccd1 _13822_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10273_ hold5210/X _10601_/B _10272_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10273_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5671 _16376_/Q vssd1 vssd1 vccd1 vccd1 hold5671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5682 _13824_/Y vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5693 _16550_/Q vssd1 vssd1 vccd1 vccd1 hold5693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ _12204_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__or2_1
Xhold4970 _16605_/Q vssd1 vssd1 vccd1 vccd1 hold4970/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4981 _10489_/X vssd1 vssd1 vccd1 vccd1 _16653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4992 _16739_/Q vssd1 vssd1 vccd1 vccd1 hold4992/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16820_ _18052_/CLK _16820_/D vssd1 vssd1 vccd1 vccd1 _16820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout470 _11594_/S vssd1 vssd1 vccd1 vccd1 _12329_/C sky130_fd_sc_hd__clkbuf_8
Xfanout481 _11480_/S vssd1 vssd1 vccd1 vccd1 _11219_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout492 _10025_/C vssd1 vssd1 vccd1 vccd1 _10019_/C sky130_fd_sc_hd__clkbuf_8
X_16751_ _17952_/CLK _16751_/D vssd1 vssd1 vccd1 vccd1 _16751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13963_ hold1408/X _13995_/A2 _13962_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _13963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15702_ _17270_/CLK _15702_/D vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ hold3383/X _12913_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16682_ _18287_/CLK _16682_/D vssd1 vssd1 vccd1 vccd1 _16682_/Q sky130_fd_sc_hd__dfxtp_1
X_13894_ _15509_/A hold1752/X hold124/X vssd1 vssd1 vccd1 vccd1 _13895_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _18421_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15633_ _17244_/CLK _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ hold3430/X _12844_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18352_ _18378_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ hold3338/X _12775_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__mux2_1
X_15564_ _17200_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17303_ _17303_/CLK _17303_/D vssd1 vssd1 vccd1 vccd1 hold830/A sky130_fd_sc_hd__dfxtp_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _14910_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14515_/X sky130_fd_sc_hd__or2_1
X_11727_ hold3563/X _11631_/A _11726_/X vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__a21oi_1
X_18283_ _18379_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ hold999/X hold1173/X hold691/X vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17234_ _17234_/CLK _17234_/D vssd1 vssd1 vccd1 vccd1 _17234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11658_ _11658_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11658_/X sky130_fd_sc_hd__or2_1
X_14446_ hold2951/X _14446_/A2 _14445_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _18461_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _16693_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_153_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14377_ hold181/X hold426/X hold333/X vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__mux2_1
X_17165_ _17198_/CLK _17165_/D vssd1 vssd1 vccd1 vccd1 _17165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11589_ _12219_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold907 hold907/A vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold918 input3/X vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ _17339_/CLK _16116_/D vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__dfxtp_1
X_13328_ hold1188/X _17563_/Q _13622_/S vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_17096_ _17160_/CLK _17096_/D vssd1 vssd1 vccd1 vccd1 _17096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _16095_/CLK _16047_/D vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__dfxtp_1
X_13259_ _13258_/X hold5920/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__mux2_1
Xhold3009 _15194_/X vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2308 _18340_/Q vssd1 vssd1 vccd1 vccd1 hold2308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2319 _17795_/Q vssd1 vssd1 vccd1 vccd1 hold2319/X sky130_fd_sc_hd__dlygate4sd3_1
X_07820_ hold531/X _14555_/C _14735_/A _09495_/C vssd1 vssd1 vccd1 vccd1 _09122_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_100_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1607 _18202_/Q vssd1 vssd1 vccd1 vccd1 hold1607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _16254_/Q vssd1 vssd1 vccd1 vccd1 hold1618/X sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _18030_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1629 _08202_/X vssd1 vssd1 vccd1 vccd1 _15737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ _18062_/CLK _16949_/D vssd1 vssd1 vccd1 vccd1 _16949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09421_ _07804_/A _09463_/B _15304_/A _09420_/X vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ hold246/A hold469/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09366_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_133_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_416_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17908_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _14862_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09283_ _15559_/A hold1517/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09283_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _14794_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08165_ _12804_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__and2_1
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08096_ _14782_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__or2_1
Xhold4200 _15283_/X vssd1 vssd1 vccd1 vccd1 _15284_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4211 _16742_/Q vssd1 vssd1 vccd1 vccd1 hold4211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4222 _11881_/X vssd1 vssd1 vccd1 vccd1 _17117_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4233 _17172_/Q vssd1 vssd1 vccd1 vccd1 hold4233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4244 _13468_/X vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3510 _13654_/X vssd1 vssd1 vccd1 vccd1 _17671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4255 _17684_/Q vssd1 vssd1 vccd1 vccd1 hold4255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3521 _17397_/Q vssd1 vssd1 vccd1 vccd1 hold3521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4266 _11638_/X vssd1 vssd1 vccd1 vccd1 _17036_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3532 _13561_/X vssd1 vssd1 vccd1 vccd1 _17640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4277 _17023_/Q vssd1 vssd1 vccd1 vccd1 hold4277/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3543 _16519_/Q vssd1 vssd1 vccd1 vccd1 hold3543/X sky130_fd_sc_hd__buf_2
Xhold4288 _13747_/X vssd1 vssd1 vccd1 vccd1 _17702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3554 _10590_/Y vssd1 vssd1 vccd1 vccd1 _10591_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4299 _16841_/Q vssd1 vssd1 vccd1 vccd1 hold4299/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2820 _15540_/X vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3565 _17562_/Q vssd1 vssd1 vccd1 vccd1 hold3565/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2831 _14619_/X vssd1 vssd1 vccd1 vccd1 _18101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3576 _10644_/Y vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08998_ _12444_/A hold479/X vssd1 vssd1 vccd1 vccd1 _16116_/D sky130_fd_sc_hd__and2_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3587 _12551_/X vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2842 _17931_/Q vssd1 vssd1 vccd1 vccd1 hold2842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2853 _14769_/X vssd1 vssd1 vccd1 vccd1 _18173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3598 _17497_/Q vssd1 vssd1 vccd1 vccd1 hold3598/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 _15703_/Q vssd1 vssd1 vccd1 vccd1 hold2864/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2875 _14442_/X vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ hold2042/X _07991_/A2 _07948_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _07949_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2886 _18058_/Q vssd1 vssd1 vccd1 vccd1 hold2886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2897 _08314_/X vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ hold3884/X _11726_/B _10959_/X _12981_/A vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09619_ hold3970/X _10007_/B _09618_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10891_ hold5304/X _11177_/B _10890_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _12789_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _17386_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_157_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17298_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12561_ _12960_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _17363_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14300_ _14910_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__or2_1
X_11512_ hold4491/X _12344_/B _11511_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11512_/X
+ sky130_fd_sc_hd__o211a_1
X_15280_ hold318/X _15486_/A2 _09357_/B _16057_/Q vssd1 vssd1 vccd1 vccd1 _15280_/X
+ sky130_fd_sc_hd__a22o_1
X_12492_ _17339_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ hold2453/X _14216_/Y _14230_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14231_/X
+ sky130_fd_sc_hd__o211a_1
X_11443_ hold4179/X _11729_/B _11442_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ _14843_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__nor2_1
X_11374_ hold5497/X _11762_/B _11373_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11374_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13113_ _13113_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__and2_1
XFILLER_0_225_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ hold1529/X _16599_/Q _10613_/C vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__mux2_1
X_14093_ hold2858/X _14094_/B _14092_/Y _14356_/A vssd1 vssd1 vccd1 vccd1 _14093_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ hold990/X hold954/X _13043_/X _13029_/A vssd1 vssd1 vccd1 vccd1 _13044_/X
+ sky130_fd_sc_hd__a211o_1
X_17921_ _18016_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5490 _12229_/X vssd1 vssd1 vccd1 vccd1 _17233_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10256_ hold1664/X hold3962/X _10997_/S vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ _17852_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10187_ hold2652/X hold3659/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16803_ _18064_/CLK _16803_/D vssd1 vssd1 vccd1 vccd1 _16803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _17975_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14995_ hold1943/X hold514/X _14994_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16734_ _17892_/CLK _16734_/D vssd1 vssd1 vccd1 vccd1 _16734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13946_ _14627_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_233_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16665_ _18221_/CLK _16665_/D vssd1 vssd1 vccd1 vccd1 _16665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13877_ _17746_/Q _13877_/B _13877_/C vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__and3_1
XFILLER_0_76_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18404_ _18404_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15616_ _17198_/CLK _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12828_ _12912_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _17452_/D sky130_fd_sc_hd__and2_1
X_16596_ _18152_/CLK _16596_/D vssd1 vssd1 vccd1 vccd1 _16596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18335_ _18341_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15547_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12759_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _17429_/D sky130_fd_sc_hd__and2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ _18266_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
X_15478_ hold431/X _09367_/A _15488_/A2 hold443/X vssd1 vssd1 vccd1 vccd1 _15478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _17217_/CLK _17217_/D vssd1 vssd1 vccd1 vccd1 _17217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14429_ _15543_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18197_ _18229_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold704 hold704/A vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ _17276_/CLK _17148_/D vssd1 vssd1 vccd1 vccd1 _17148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold715 hold715/A vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 hold726/A vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 hold737/A vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ hold5206/X _10571_/B _09969_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _09970_/X
+ sky130_fd_sc_hd__o211a_1
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _17970_/CLK _17079_/D vssd1 vssd1 vccd1 vccd1 _17079_/Q sky130_fd_sc_hd__dfxtp_1
X_08921_ _15264_/A hold223/X vssd1 vssd1 vccd1 vccd1 _16078_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2105 _13989_/X vssd1 vssd1 vccd1 vccd1 _17799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 _14825_/X vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08852_ hold578/X hold615/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__mux2_1
Xhold2127 _12975_/X vssd1 vssd1 vccd1 vccd1 _17501_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2138 _16208_/Q vssd1 vssd1 vccd1 vccd1 hold2138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 _17513_/Q vssd1 vssd1 vccd1 vccd1 hold1404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _15659_/Q vssd1 vssd1 vccd1 vccd1 hold2149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _08218_/X vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07803_ _16286_/Q _07801_/B _07802_/Y vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__o21ai_1
Xhold1426 _07935_/X vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ hold210/X _16012_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__mux2_1
Xhold1437 _07880_/X vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1448 _17895_/Q vssd1 vssd1 vccd1 vccd1 hold1448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _14331_/X vssd1 vssd1 vccd1 vccd1 _17963_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09404_ _09438_/B _09404_/B vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_250_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18166_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09335_ _15231_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _12747_/A hold447/X vssd1 vssd1 vccd1 vccd1 hold448/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08217_ _14330_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__or2_1
X_09197_ hold3049/X _09218_/B _09196_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _09197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08148_ _14726_/A hold2522/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_6_44_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_44_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_08079_ hold2471/X _08088_/B _08078_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08079_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4030 _16970_/Q vssd1 vssd1 vccd1 vccd1 hold4030/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4041 _09925_/X vssd1 vssd1 vccd1 vccd1 _16465_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10110_ _10554_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__or2_1
XTAP_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4052 _17723_/Q vssd1 vssd1 vccd1 vccd1 hold4052/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4063 _16493_/Q vssd1 vssd1 vccd1 vccd1 hold4063/X sky130_fd_sc_hd__dlygate4sd3_1
X_11090_ hold3213/X _16854_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _11091_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4074 _13525_/X vssd1 vssd1 vccd1 vccd1 _17628_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4085 _17154_/Q vssd1 vssd1 vccd1 vccd1 hold4085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3340 _17387_/Q vssd1 vssd1 vccd1 vccd1 hold3340/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3351 _16456_/Q vssd1 vssd1 vccd1 vccd1 hold3351/X sky130_fd_sc_hd__dlygate4sd3_1
X_10041_ _13222_/A _10191_/A _10040_/X vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__a21oi_1
Xhold4096 _10993_/X vssd1 vssd1 vccd1 vccd1 _16821_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3362 _09517_/X vssd1 vssd1 vccd1 vccd1 _16329_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3373 _12722_/X vssd1 vssd1 vccd1 vccd1 _12723_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__buf_6
Xhold3384 _16359_/Q vssd1 vssd1 vccd1 vccd1 hold3384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3395 _17693_/Q vssd1 vssd1 vccd1 vccd1 hold3395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2650 _15772_/Q vssd1 vssd1 vccd1 vccd1 hold2650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__buf_4
XFILLER_0_227_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2661 _08292_/X vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2672 _15856_/Q vssd1 vssd1 vccd1 vccd1 hold2672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 _17892_/Q vssd1 vssd1 vccd1 vccd1 hold2683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 _14548_/X vssd1 vssd1 vccd1 vccd1 _18068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1960 _18070_/Q vssd1 vssd1 vccd1 vccd1 hold1960/X sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _13800_/A _13800_/B vssd1 vssd1 vccd1 vccd1 _13800_/X sky130_fd_sc_hd__or2_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_338_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17215_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1971 _14881_/X vssd1 vssd1 vccd1 vccd1 _18227_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14780_ _15227_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__or2_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11992_ hold4153/X _12374_/B _11991_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11992_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1982 _14951_/X vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1993 _08192_/X vssd1 vssd1 vccd1 vccd1 _15732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10943_ hold3041/X hold5487/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__mux2_1
X_13731_ _13767_/A _13731_/B vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16450_ _18265_/CLK _16450_/D vssd1 vssd1 vccd1 vccd1 _16450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ hold2545/X _16782_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13662_ _13788_/A _13662_/B vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15401_ _16304_/Q _09362_/A _09392_/B hold876/X _15400_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/D sky130_fd_sc_hd__a221o_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12613_ hold1432/X _17382_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16381_ _18292_/CLK _16381_/D vssd1 vssd1 vccd1 vccd1 _16381_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13593_ _13791_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18152_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15332_ _15489_/A _15332_/B _15332_/C _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_171_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12544_ hold2901/X _17359_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18051_ _18061_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ hold118/X _12445_/A _08868_/X _12474_/X _09055_/A vssd1 vssd1 vccd1 vccd1
+ hold39/A sky130_fd_sc_hd__o311a_1
X_15263_ _15490_/A1 _15255_/X _15262_/X _15490_/B1 _18400_/Q vssd1 vssd1 vccd1 vccd1
+ _15263_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ _17880_/CLK _17002_/D vssd1 vssd1 vccd1 vccd1 _17002_/Q sky130_fd_sc_hd__dfxtp_1
X_14214_ _15559_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__or2_1
X_11426_ hold1208/X hold3762/X _11711_/S vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__mux2_1
XANTENNA_6 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15194_ hold3008/X _15221_/B _15193_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _15194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18049_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14145_ hold2023/X _14148_/B _14144_/Y _13905_/A vssd1 vssd1 vccd1 vccd1 _14145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11357_ hold2961/X _16943_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11358_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10308_ _10524_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__or2_1
X_14076_ _15203_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14076_/X sky130_fd_sc_hd__or2_1
X_11288_ hold1349/X hold5004/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13027_ _13034_/D hold957/A vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__and2_1
XFILLER_0_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17904_ _17904_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_1
X_10239_ _10554_/A _10239_/B vssd1 vssd1 vccd1 vccd1 _10239_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17835_ _17867_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17766_ _17894_/CLK _17766_/D vssd1 vssd1 vccd1 vccd1 _17766_/Q sky130_fd_sc_hd__dfxtp_1
X_14978_ hold525/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16717_ _18046_/CLK _16717_/D vssd1 vssd1 vccd1 vccd1 _16717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13929_ _13929_/A hold247/X vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__and2_1
XFILLER_0_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17697_ _17729_/CLK _17697_/D vssd1 vssd1 vccd1 vccd1 _17697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16648_ _18210_/CLK _16648_/D vssd1 vssd1 vccd1 vccd1 _16648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ _18216_/CLK _16579_/D vssd1 vssd1 vccd1 vccd1 _16579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _18457_/Q _11158_/A _18460_/Q vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nor3_1
X_18318_ _18318_/CLK hold624/X vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09051_ _09055_/A hold490/X vssd1 vssd1 vccd1 vccd1 _16142_/D sky130_fd_sc_hd__and2_1
XFILLER_0_199_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _18383_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ hold2459/X _08033_/B _08001_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _08002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold501 hold558/X vssd1 vssd1 vccd1 vccd1 hold559/A sky130_fd_sc_hd__buf_6
XFILLER_0_130_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold512 hold753/X vssd1 vssd1 vccd1 vccd1 hold754/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold523 hold523/A vssd1 vssd1 vccd1 vccd1 input64/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 hold545/A vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 hold556/A vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold567 input14/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold578 hold59/X vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__buf_4
XFILLER_0_229_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ hold1851/X hold3655/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__mux2_1
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_08904_ hold379/X _16070_/Q _08928_/S vssd1 vssd1 vccd1 vccd1 hold380/A sky130_fd_sc_hd__mux2_1
XFILLER_0_209_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ hold962/X hold4026/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _18015_/Q vssd1 vssd1 vccd1 vccd1 hold1201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _18388_/Q vssd1 vssd1 vccd1 vccd1 hold1212/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _12438_/A hold435/X vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1223 _15829_/Q vssd1 vssd1 vccd1 vccd1 hold1223/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 _17777_/Q vssd1 vssd1 vccd1 vccd1 hold1234/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1245 _15828_/Q vssd1 vssd1 vccd1 vccd1 hold1245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1256 _15588_/Q vssd1 vssd1 vccd1 vccd1 hold1256/X sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ _15344_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _16003_/D sky130_fd_sc_hd__and2_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_431_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17613_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1267 _18005_/Q vssd1 vssd1 vccd1 vccd1 hold1267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _08475_/X vssd1 vssd1 vccd1 vccd1 _15866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 _15878_/Q vssd1 vssd1 vccd1 vccd1 hold1289/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08697_ hold256/X hold404/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08698_/B sky130_fd_sc_hd__mux2_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09318_ hold2933/X _09325_/B _09317_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ hold3553/X _10554_/A _10589_/X vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ _15525_/A hold3035/X _09273_/S vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ hold2669/X _17244_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ hold4929/X _11667_/A _11210_/X vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12191_ hold2441/X _17221_/Q _12302_/C vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11142_ hold3732/X _11052_/A _11141_/X vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_222_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput76 _13161_/A vssd1 vssd1 vccd1 vccd1 output76/X sky130_fd_sc_hd__buf_6
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 _13241_/A vssd1 vssd1 vccd1 vccd1 output87/X sky130_fd_sc_hd__buf_6
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _17297_/CLK _15950_/D vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__dfxtp_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073_ _11553_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__or2_1
Xoutput98 _13089_/A vssd1 vssd1 vccd1 vccd1 output98/X sky130_fd_sc_hd__buf_6
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3170 _17369_/Q vssd1 vssd1 vccd1 vccd1 hold3170/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ hold1389/X _14896_/Y _14900_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _14901_/X
+ sky130_fd_sc_hd__o211a_1
X_10024_ _11158_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _16498_/D sky130_fd_sc_hd__nor2_1
Xhold3181 _17448_/Q vssd1 vssd1 vccd1 vccd1 hold3181/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3192 _14987_/X vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _17719_/CLK _15881_/D vssd1 vssd1 vccd1 vccd1 _15881_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2480 _18241_/Q vssd1 vssd1 vccd1 vccd1 hold2480/X sky130_fd_sc_hd__dlygate4sd3_1
X_17620_ _17748_/CLK _17620_/D vssd1 vssd1 vccd1 vccd1 _17620_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2491 _14947_/X vssd1 vssd1 vccd1 vccd1 _18258_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14832_ _15225_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14832_/X sky130_fd_sc_hd__or2_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_172_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18377_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_231_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17551_ _18221_/CLK _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18411_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1790 _14631_/X vssd1 vssd1 vccd1 vccd1 _18106_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14763_ hold1931/X _14774_/B _14762_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14763_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ hold1186/X _17149_/Q _12251_/S vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__mux2_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16502_ _18323_/CLK _16502_/D vssd1 vssd1 vccd1 vccd1 _16502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13714_ _13808_/A _13802_/B _13713_/X _13714_/C1 vssd1 vssd1 vccd1 vccd1 _17691_/D
+ sky130_fd_sc_hd__o211a_1
X_10926_ _11103_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__or2_1
X_17482_ _17482_/CLK _17482_/D vssd1 vssd1 vccd1 vccd1 _17482_/Q sky130_fd_sc_hd__dfxtp_1
X_14694_ _14910_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16433_ _18386_/CLK _16433_/D vssd1 vssd1 vccd1 vccd1 _16433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10857_ _11052_/A _10857_/B vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__or2_1
X_13645_ hold4563/X _13856_/B _13644_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13645_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _18309_/CLK _16364_/D vssd1 vssd1 vccd1 vccd1 _16364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ hold5719/X _13829_/B _13575_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13576_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _11070_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18216_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_1
X_15315_ hold727/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ hold3261/X _12526_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16295_ _16323_/CLK _16295_/D vssd1 vssd1 vccd1 vccd1 _16295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18034_ _18068_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _17328_/Q _15448_/B1 _15485_/B1 hold457/X vssd1 vssd1 vccd1 vccd1 _15246_/X
+ sky130_fd_sc_hd__a22o_1
X_12458_ _17322_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_239_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11409_ _12246_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ _15231_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__or2_1
X_12389_ hold88/X hold129/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ _14862_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ hold1359/X _14107_/A2 _14058_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _14059_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08620_ _09015_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _15932_/D sky130_fd_sc_hd__and2_1
XFILLER_0_193_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17818_ _17822_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _12418_/A hold707/X vssd1 vssd1 vccd1 vccd1 _15899_/D sky130_fd_sc_hd__and2_1
X_17749_ _17749_/CLK _17749_/D vssd1 vssd1 vccd1 vccd1 _17749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08482_ _15541_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09103_ hold2025/X _09106_/B _09102_/Y _12975_/A vssd1 vssd1 vccd1 vccd1 _09103_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ hold379/X hold616/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__buf_2
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold342 hold342/A vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold56/X vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__buf_4
Xhold364 la_data_in[19] vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/A vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 hold386/A vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout800 _15068_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__buf_4
Xhold397 hold397/A vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _15192_/C1 vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__buf_4
XFILLER_0_217_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__or2_1
Xfanout822 _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14813_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout833 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14883_/C1 sky130_fd_sc_hd__buf_2
Xfanout844 _14815_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/C1 sky130_fd_sc_hd__buf_4
Xfanout855 _15004_/A vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__buf_12
XFILLER_0_42_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout866 fanout873/X vssd1 vssd1 vccd1 vccd1 _12367_/A sky130_fd_sc_hd__buf_6
XFILLER_0_102_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09867_ _09963_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09867_/X sky130_fd_sc_hd__or2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 hold943/X vssd1 vssd1 vccd1 vccd1 hold944/A sky130_fd_sc_hd__clkbuf_2
Xfanout888 hold525/X vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__clkbuf_16
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 hold1020/A vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__clkbuf_16
Xhold1031 _15141_/X vssd1 vssd1 vccd1 vccd1 hold1031/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout899 _14972_/A vssd1 vssd1 vccd1 vccd1 _15513_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1042 _17977_/Q vssd1 vssd1 vccd1 vccd1 hold1042/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ hold596/X hold786/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold787/A sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1053 _09183_/X vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _09936_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__or2_1
Xhold1064 _09079_/X vssd1 vssd1 vccd1 vccd1 _16154_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1075 _15088_/X vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _08425_/X vssd1 vssd1 vccd1 vccd1 hold1086/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _08233_/X vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08749_ hold163/X _15995_/Q _08779_/S vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ hold5102/X _11670_/A _11759_/X vssd1 vssd1 vccd1 vccd1 _11760_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_240_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ hold5078/X _11095_/A2 _10710_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _10711_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _12234_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ _11218_/A _10642_/B vssd1 vssd1 vccd1 vccd1 _16704_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13430_ hold2174/X _17597_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ hold2195/X hold3702/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ _10603_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _16681_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ hold2963/X _15113_/B _15099_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _15100_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12312_ hold4787/X _12261_/A _12311_/X vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16080_ _18399_/CLK _16080_/D vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13292_ hold3850/X _13291_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13292_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15031_ _15193_/A hold2544/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15032_/B sky130_fd_sc_hd__mux2_1
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ _12273_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ hold4537/X _11207_/B _11124_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11125_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_353_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17740_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16982_ _17935_/CLK _16982_/D vssd1 vssd1 vccd1 vccd1 _16982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15933_ _16097_/CLK _15933_/D vssd1 vssd1 vccd1 vccd1 hold431/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ hold3401/X _11150_/B _11055_/X _12981_/A vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _16493_/Q _10007_/B _10007_/C vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__and3_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _17217_/CLK _15864_/D vssd1 vssd1 vccd1 vccd1 _15864_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _17667_/CLK _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
X_14815_ hold2935/X _14826_/B _14814_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _14815_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _17726_/CLK _15795_/D vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17534_/CLK _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14746_ _15193_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14746_/X sky130_fd_sc_hd__or2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11958_ _12246_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10909_ hold4240/X _11180_/B _10908_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17465_ _17483_/CLK _17465_/D vssd1 vssd1 vccd1 vccd1 _17465_/Q sky130_fd_sc_hd__dfxtp_1
X_14677_ hold1509/X _14664_/B _14676_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ _12273_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16416_ _18327_/CLK _16416_/D vssd1 vssd1 vccd1 vccd1 _16416_/Q sky130_fd_sc_hd__dfxtp_1
X_13628_ hold2047/X hold5707/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17396_ _18445_/CLK _17396_/D vssd1 vssd1 vccd1 vccd1 _17396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ _18360_/CLK _16347_/D vssd1 vssd1 vccd1 vccd1 _16347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ hold2194/X _17640_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6009 data_in[31] vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _17510_/CLK _16278_/D vssd1 vssd1 vccd1 vccd1 _16278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5308 _17235_/Q vssd1 vssd1 vccd1 vccd1 hold5308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5319 _11008_/X vssd1 vssd1 vccd1 vccd1 _16826_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18017_ _18017_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
X_15229_ _15229_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4607 _10575_/Y vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4618 _10650_/Y vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4629 _16340_/Q vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3906 _16681_/Q vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3917 _10456_/X vssd1 vssd1 vccd1 vccd1 _16642_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3928 _16936_/Q vssd1 vssd1 vccd1 vccd1 hold3928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3939 _13510_/X vssd1 vssd1 vccd1 vccd1 _17623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07982_ _15551_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07982_/X sky130_fd_sc_hd__or2_1
X_09721_ hold4137/X _10007_/B _09720_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09721_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ hold3365/X _10004_/B _09651_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09652_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08603_ hold215/X hold759/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__mux2_1
X_09583_ hold4713/X _10577_/B _09582_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ hold312/X hold506/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold507/A sky130_fd_sc_hd__mux2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08465_ hold1630/X _08488_/B _08464_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _08465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ hold1245/X _08440_/A2 _08395_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ _09055_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _16125_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5820 hold5947/X vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__buf_1
XFILLER_0_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5831 _18404_/Q vssd1 vssd1 vccd1 vccd1 hold5831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5842 hold5842/A vssd1 vssd1 vccd1 vccd1 hold5842/X sky130_fd_sc_hd__buf_2
Xhold5853 _18399_/Q vssd1 vssd1 vccd1 vccd1 hold5853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hold8/X vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__buf_4
Xhold5864 hold5864/A vssd1 vssd1 vccd1 vccd1 hold5864/X sky130_fd_sc_hd__clkbuf_4
Xhold5875 _18419_/Q vssd1 vssd1 vccd1 vccd1 hold5875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 hold64/X vssd1 vssd1 vccd1 vccd1 input36/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5886 hold5886/A vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_12
Xhold172 hold25/X vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5897 _17752_/Q vssd1 vssd1 vccd1 vccd1 hold5897/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout630 _09440_/X vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__clkbuf_4
Xfanout641 _12807_/A vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__buf_4
X_09919_ hold3379/X _10013_/B _09918_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout652 _12909_/A vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__buf_4
Xfanout663 _12981_/A vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout674 _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__buf_2
Xfanout685 fanout692/X vssd1 vssd1 vccd1 vccd1 _14554_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_226_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout696 _12600_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__buf_4
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _12996_/A _12930_/B vssd1 vssd1 vccd1 vccd1 _17486_/D sky130_fd_sc_hd__and2_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12861_ _12870_/A _12861_/B vssd1 vssd1 vccd1 vccd1 _17463_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14600_ _15209_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__or2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ hold5232/X _13798_/A2 _11811_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11812_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _17280_/CLK _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12807_/A _12792_/B vssd1 vssd1 vccd1 vccd1 _17440_/D sky130_fd_sc_hd__and2_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _15103_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__or2_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13864_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _17071_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17250_ _17607_/CLK _17250_/D vssd1 vssd1 vccd1 vccd1 _17250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ hold2733/X _14482_/A2 _14461_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14462_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ hold5629/X _11768_/B _11673_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11674_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16201_ _17507_/CLK _16201_/D vssd1 vssd1 vccd1 vccd1 _16201_/Q sky130_fd_sc_hd__dfxtp_1
X_13413_ _13797_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ _16699_/Q _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__and3_1
XFILLER_0_183_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17181_ _17245_/CLK _17181_/D vssd1 vssd1 vccd1 vccd1 _17181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_3_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ hold733/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _17327_/CLK _16132_/D vssd1 vssd1 vccd1 vccd1 _16132_/Q sky130_fd_sc_hd__dfxtp_1
X_10556_ hold1214/X hold3643/X _11096_/S vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__mux2_1
X_13344_ _13767_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _18408_/CLK _16063_/D vssd1 vssd1 vccd1 vccd1 hold847/A sky130_fd_sc_hd__dfxtp_1
X_10487_ hold1933/X hold4968/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10488_/B sky130_fd_sc_hd__mux2_1
X_13275_ _13274_/X hold4998/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15014_ _15121_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12226_ hold5340/X _12353_/B _12225_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ hold3432/X _12347_/B _12156_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ hold2909/X hold4427/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12088_ hold4143/X _12374_/B _12087_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__o211a_1
X_16965_ _17875_/CLK _16965_/D vssd1 vssd1 vccd1 vccd1 _16965_/Q sky130_fd_sc_hd__dfxtp_1
X_15916_ _16322_/CLK _15916_/D vssd1 vssd1 vccd1 vccd1 hold679/A sky130_fd_sc_hd__dfxtp_1
X_11039_ hold2937/X hold5543/X _11156_/C vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_223_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16896_ _18065_/CLK _16896_/D vssd1 vssd1 vccd1 vccd1 _16896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _17703_/CLK _15847_/D vssd1 vssd1 vccd1 vccd1 _15847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _17613_/CLK _15778_/D vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfxtp_1
X_17517_ _17517_/CLK _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_1
X_14729_ hold2339/X _14720_/B _14728_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ _15203_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _17455_/CLK _17448_/D vssd1 vssd1 vccd1 vccd1 _17448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ _15515_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__or2_1
X_17379_ _17379_/CLK _17379_/D vssd1 vssd1 vccd1 vccd1 _17379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5105 _09724_/X vssd1 vssd1 vccd1 vccd1 _16398_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5116 _17137_/Q vssd1 vssd1 vccd1 vccd1 hold5116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5127 _10474_/X vssd1 vssd1 vccd1 vccd1 _16648_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_275_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18170_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5138 _17598_/Q vssd1 vssd1 vccd1 vccd1 hold5138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5149 _10720_/X vssd1 vssd1 vccd1 vccd1 _16730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4404 _10717_/X vssd1 vssd1 vccd1 vccd1 _16729_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4415 _16872_/Q vssd1 vssd1 vccd1 vccd1 hold4415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4426 _10921_/X vssd1 vssd1 vccd1 vccd1 _16797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_204_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18292_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4437 _17056_/Q vssd1 vssd1 vccd1 vccd1 hold4437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4448 _15433_/X vssd1 vssd1 vccd1 vccd1 _15434_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3703 _13842_/Y vssd1 vssd1 vccd1 vccd1 _13843_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3714 _16688_/Q vssd1 vssd1 vccd1 vccd1 hold3714/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4459 _16862_/Q vssd1 vssd1 vccd1 vccd1 hold4459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3725 _12342_/Y vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3736 _17121_/Q vssd1 vssd1 vccd1 vccd1 hold3736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3747 _11521_/X vssd1 vssd1 vccd1 vccd1 _16997_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3758 _16713_/Q vssd1 vssd1 vccd1 vccd1 hold3758/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3769 _09799_/X vssd1 vssd1 vccd1 vccd1 _16423_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07965_ hold2743/X _07978_/B _07964_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _07965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09704_ hold1005/X hold3966/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07896_ _14854_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ hold2995/X _16369_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09566_ hold1491/X _13238_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08517_ _15521_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _15551_/A _15169_/A hold246/A _15215_/A vssd1 vssd1 vccd1 vccd1 _09498_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08448_ hold202/X _14913_/A vssd1 vssd1 vccd1 vccd1 _08448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08379_ _08379_/A hold664/X vssd1 vssd1 vccd1 vccd1 _15821_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10410_ _10542_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11390_ hold1265/X _16954_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10341_ _10497_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ hold4155/X _13059_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
Xhold5650 _17045_/Q vssd1 vssd1 vccd1 vccd1 hold5650/X sky130_fd_sc_hd__dlygate4sd3_1
X_10272_ _10488_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__or2_1
Xhold5661 _16380_/Q vssd1 vssd1 vccd1 vccd1 hold5661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5672 _09562_/X vssd1 vssd1 vccd1 vccd1 _16344_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5683 _16418_/Q vssd1 vssd1 vccd1 vccd1 hold5683/X sky130_fd_sc_hd__dlygate4sd3_1
X_12011_ hold2785/X _17161_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5694 _10084_/X vssd1 vssd1 vccd1 vccd1 _16518_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4960 _16731_/Q vssd1 vssd1 vccd1 vccd1 hold4960/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4971 _10249_/X vssd1 vssd1 vccd1 vccd1 _16573_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4982 _17051_/Q vssd1 vssd1 vccd1 vccd1 hold4982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4993 _11226_/Y vssd1 vssd1 vccd1 vccd1 _11227_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout460 _10025_/C vssd1 vssd1 vccd1 vccd1 _13847_/C sky130_fd_sc_hd__buf_4
XFILLER_0_217_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout471 _11594_/S vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__clkbuf_8
X_16750_ _18060_/CLK _16750_/D vssd1 vssd1 vccd1 vccd1 _16750_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout482 _10025_/C vssd1 vssd1 vccd1 vccd1 _11480_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout493 _10001_/C vssd1 vssd1 vccd1 vccd1 _10007_/C sky130_fd_sc_hd__clkbuf_8
X_13962_ _15523_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15701_ _17237_/CLK _15701_/D vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_79_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17370_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ hold2768/X hold3315/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_220_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16681_ _18233_/CLK _16681_/D vssd1 vssd1 vccd1 vccd1 _16681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13893_ hold238/X hold122/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__nand2_1
XFILLER_0_198_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18420_ _18422_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_159_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15632_ _17157_/CLK _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ hold1881/X hold3419/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_201_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18351_ _18351_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15563_ _17263_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ hold2562/X _17436_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17303_/CLK _17302_/D vssd1 vssd1 vccd1 vccd1 hold792/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14514_ hold2892/X _14535_/B _14513_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14514_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18380_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _17066_/Q _11726_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15494_ _15494_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17233_ _17900_/CLK _17233_/D vssd1 vssd1 vccd1 vccd1 _17233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ _15233_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14445_/X sky130_fd_sc_hd__or2_1
X_11657_ hold2329/X hold5529/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ hold4637/X _10536_/A _10607_/X vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__a21oi_1
X_17164_ _17164_/CLK _17164_/D vssd1 vssd1 vccd1 vccd1 _17164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14376_ _14376_/A hold334/X vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__and2_1
X_11588_ hold2345/X hold5124/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16115_ _17343_/CLK _16115_/D vssd1 vssd1 vccd1 vccd1 _16115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold908 hold908/A vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ hold3942/X _13802_/B _13326_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13327_/X
+ sky130_fd_sc_hd__o211a_1
Xhold919 hold953/X vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ _11100_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17095_ _17221_/CLK _17095_/D vssd1 vssd1 vccd1 vccd1 _17095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ _16127_/CLK _16046_/D vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13258_ _17583_/Q _17117_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13258_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ hold1425/X _17227_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13188_/X hold4630/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13189_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2309 _15116_/X vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1608 _14829_/X vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _17997_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1619 _09288_/X vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16948_ _17858_/CLK _16948_/D vssd1 vssd1 vccd1 vccd1 _16948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16879_ _17952_/CLK _16879_/D vssd1 vssd1 vccd1 vccd1 _16879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ _09438_/B _16296_/Q vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09351_ _09366_/A _09351_/B _09360_/B vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08302_ hold1979/X _08336_/A2 _08301_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08302_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09282_ _12696_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _16252_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08233_ hold1096/X _08263_/A2 _08232_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_456_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17689_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _15515_/A hold2526/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08095_ hold2741/X _08097_/A2 _08094_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _08095_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_34_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_34_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4201 _17199_/Q vssd1 vssd1 vccd1 vccd1 hold4201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4212 _10660_/X vssd1 vssd1 vccd1 vccd1 _16710_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4223 _16806_/Q vssd1 vssd1 vccd1 vccd1 hold4223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4234 _11950_/X vssd1 vssd1 vccd1 vccd1 _17140_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3500 _17745_/Q vssd1 vssd1 vccd1 vccd1 hold3500/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4245 _17748_/Q vssd1 vssd1 vccd1 vccd1 hold4245/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4256 _13597_/X vssd1 vssd1 vccd1 vccd1 _17652_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3511 _17711_/Q vssd1 vssd1 vccd1 vccd1 hold3511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3522 _12662_/X vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4267 _17246_/Q vssd1 vssd1 vccd1 vccd1 hold4267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3533 _16875_/Q vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4278 _11503_/X vssd1 vssd1 vccd1 vccd1 _16991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3544 _10566_/Y vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4289 _17251_/Q vssd1 vssd1 vccd1 vccd1 hold4289/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3555 _16538_/Q vssd1 vssd1 vccd1 vccd1 hold3555/X sky130_fd_sc_hd__buf_1
Xhold2810 _18065_/Q vssd1 vssd1 vccd1 vccd1 hold2810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3566 _13806_/Y vssd1 vssd1 vccd1 vccd1 _13807_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2821 _17819_/Q vssd1 vssd1 vccd1 vccd1 hold2821/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3577 _17379_/Q vssd1 vssd1 vccd1 vccd1 hold3577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 _16199_/Q vssd1 vssd1 vccd1 vccd1 hold2832/X sky130_fd_sc_hd__dlygate4sd3_1
X_08997_ hold150/X hold478/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold479/A sky130_fd_sc_hd__mux2_1
XFILLER_0_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2843 _14265_/X vssd1 vssd1 vccd1 vccd1 _17931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3588 _17359_/Q vssd1 vssd1 vccd1 vccd1 hold3588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3599 _17364_/Q vssd1 vssd1 vccd1 vccd1 hold3599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2854 _17815_/Q vssd1 vssd1 vccd1 vccd1 hold2854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2865 _18182_/Q vssd1 vssd1 vccd1 vccd1 hold2865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2876 _16277_/Q vssd1 vssd1 vccd1 vccd1 hold2876/X sky130_fd_sc_hd__dlygate4sd3_1
X_07948_ _14403_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07948_/X sky130_fd_sc_hd__or2_1
Xhold2887 _14528_/X vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2898 _18306_/Q vssd1 vssd1 vccd1 vccd1 hold2898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07879_ _15557_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _09936_/A _09618_/B vssd1 vssd1 vccd1 vccd1 _09618_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _11082_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _09954_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ hold3606/X _12559_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _12057_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_197_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18316_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ hold32/X _12509_/A2 _12507_/A3 _12490_/X _09015_/A vssd1 vssd1 vccd1 vccd1
+ hold33/A sky130_fd_sc_hd__o311a_1
XFILLER_0_62_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _15521_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14230_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17314_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _11637_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ _11667_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__or2_1
X_14161_ hold864/X _14148_/B _14160_/X _15496_/A vssd1 vssd1 vccd1 vccd1 hold865/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13112_ _13105_/X _13111_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17532_/D sky130_fd_sc_hd__o21a_1
X_10324_ hold4022/X _10628_/B _10323_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _15545_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5480 _10846_/X vssd1 vssd1 vccd1 vccd1 _16772_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13043_ _17523_/Q hold960/X _13043_/C vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__or3_1
X_10255_ hold3726/X _10631_/B _10254_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5491 _16812_/Q vssd1 vssd1 vccd1 vccd1 hold5491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _17952_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4790 _10156_/X vssd1 vssd1 vccd1 vccd1 _16542_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17851_ _17851_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_1
X_10186_ hold4799/X _10571_/B _10185_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16802_ _18035_/CLK _16802_/D vssd1 vssd1 vccd1 vccd1 _16802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _17814_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14994_ _15209_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__or2_1
Xfanout290 _11679_/A vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__buf_2
XFILLER_0_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16733_ _17966_/CLK _16733_/D vssd1 vssd1 vccd1 vccd1 _16733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13945_ _15494_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _17778_/D sky130_fd_sc_hd__and2_1
XFILLER_0_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16664_ _17968_/CLK _16664_/D vssd1 vssd1 vccd1 vccd1 _16664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _13888_/A _13876_/B vssd1 vssd1 vccd1 vccd1 _17745_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_232_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18403_ _18403_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_2
X_15615_ _17179_/CLK _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12827_ hold3179/X _12826_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16595_ _18175_/CLK _16595_/D vssd1 vssd1 vccd1 vccd1 _16595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _18366_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ hold2518/X _15547_/B _15545_/Y _15548_/C1 vssd1 vssd1 vccd1 vccd1 _15546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ hold3674/X _12757_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18265_ _18265_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _12285_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__or2_1
X_15477_ _07805_/A _15477_/A2 _09365_/B hold767/X vssd1 vssd1 vccd1 vccd1 _15480_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ hold4139/X _12688_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17216_ _17280_/CLK _17216_/D vssd1 vssd1 vccd1 vccd1 _17216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ hold2570/X _14433_/B _14427_/Y _14362_/A vssd1 vssd1 vccd1 vccd1 _14428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18196_ _18228_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17147_ _17179_/CLK _17147_/D vssd1 vssd1 vccd1 vccd1 _17147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold705 hold705/A vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ hold944/X hold1042/X hold333/X vssd1 vssd1 vccd1 vccd1 _14360_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold716 hold716/A vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold738 hold738/A vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold749 la_data_in[26] vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
X_17078_ _17935_/CLK _17078_/D vssd1 vssd1 vccd1 vccd1 _17078_/Q sky130_fd_sc_hd__dfxtp_1
X_16029_ _17301_/CLK _16029_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
X_08920_ hold222/X _16078_/Q _08928_/S vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2106 _15695_/Q vssd1 vssd1 vccd1 vccd1 hold2106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2117 _15714_/Q vssd1 vssd1 vccd1 vccd1 hold2117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08851_ _12418_/A hold738/X vssd1 vssd1 vccd1 vccd1 _16044_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2128 _15845_/Q vssd1 vssd1 vccd1 vccd1 hold2128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2139 _09193_/X vssd1 vssd1 vccd1 vccd1 _16208_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1405 _13010_/X vssd1 vssd1 vccd1 vccd1 _17513_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ _09339_/B _07802_/B vssd1 vssd1 vccd1 vccd1 _07802_/Y sky130_fd_sc_hd__nand2_1
Xhold1416 _18047_/Q vssd1 vssd1 vccd1 vccd1 hold1416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _15594_/Q vssd1 vssd1 vccd1 vccd1 hold1427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08782_ _15454_/A hold386/X vssd1 vssd1 vccd1 vccd1 _16011_/D sky130_fd_sc_hd__and2_1
Xhold1438 la_data_in[3] vssd1 vssd1 vccd1 vccd1 hold1438/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1449 _14189_/X vssd1 vssd1 vccd1 vccd1 _17895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09403_ _07785_/Y _07786_/A _11158_/A vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09334_ hold2876/X _09338_/A2 _09333_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_290_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09265_ hold469/A _16244_/Q _09273_/S vssd1 vssd1 vccd1 vccd1 hold447/A sky130_fd_sc_hd__mux2_1
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ hold2359/X _08213_/B _08215_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09196_ _15525_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ _15537_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__or2_1
Xhold4020 _16390_/Q vssd1 vssd1 vccd1 vccd1 hold4020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4031 _11344_/X vssd1 vssd1 vccd1 vccd1 _16938_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4042 _16578_/Q vssd1 vssd1 vccd1 vccd1 hold4042/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4053 _16662_/Q vssd1 vssd1 vccd1 vccd1 hold4053/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4064 _09913_/X vssd1 vssd1 vccd1 vccd1 _16461_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4075 _16706_/Q vssd1 vssd1 vccd1 vccd1 hold4075/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3330 _17446_/Q vssd1 vssd1 vccd1 vccd1 hold3330/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _16504_/Q _10070_/B _10190_/S vssd1 vssd1 vccd1 vccd1 _10040_/X sky130_fd_sc_hd__and3_1
Xhold4086 _11896_/X vssd1 vssd1 vccd1 vccd1 _17122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3341 _17386_/Q vssd1 vssd1 vccd1 vccd1 hold3341/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3352 _09802_/X vssd1 vssd1 vccd1 vccd1 _16424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4097 _16420_/Q vssd1 vssd1 vccd1 vccd1 hold4097/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3363 _16488_/Q vssd1 vssd1 vccd1 vccd1 hold3363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3374 _16325_/Q vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__buf_4
Xhold3385 _09511_/X vssd1 vssd1 vccd1 vccd1 _16327_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 _15627_/Q vssd1 vssd1 vccd1 vccd1 hold2640/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3396 _13624_/X vssd1 vssd1 vccd1 vccd1 _17661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2651 _08275_/X vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2662 _16240_/Q vssd1 vssd1 vccd1 vccd1 hold2662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkbuf_2
Xhold2673 _08455_/X vssd1 vssd1 vccd1 vccd1 _15856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2684 _14183_/X vssd1 vssd1 vccd1 vccd1 _17892_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 _18097_/Q vssd1 vssd1 vccd1 vccd1 hold1950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2695 _18395_/Q vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 _14552_/X vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__buf_4
XFILLER_0_199_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _13461_/A _11991_/B vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__or2_1
Xhold1972 _18427_/Q vssd1 vssd1 vccd1 vccd1 hold1972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 _18380_/Q vssd1 vssd1 vccd1 vccd1 hold1983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1994 _18250_/Q vssd1 vssd1 vccd1 vccd1 hold1994/X sky130_fd_sc_hd__dlygate4sd3_1
X_13730_ hold2575/X _17697_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13731_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10942_ hold4119/X _11729_/B _10941_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _10942_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_378_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17667_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13661_ hold1706/X _17674_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10873_ hold5264/X _11159_/B _10872_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _10873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15400_ hold628/X _09367_/A _09357_/B hold442/X vssd1 vssd1 vccd1 vccd1 _15400_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ _13002_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _17380_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16380_ _18323_/CLK _16380_/D vssd1 vssd1 vccd1 vccd1 _16380_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_307_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17894_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13592_ hold1979/X _17651_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__mux2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15331_ _16297_/Q _15477_/A2 _15487_/B1 hold639/X _15330_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/D sky130_fd_sc_hd__a221o_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12606_/A _12543_/B vssd1 vssd1 vccd1 vccd1 _17357_/D sky130_fd_sc_hd__and2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _18050_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ _15489_/A _15262_/B _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _17330_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17001_ _17880_/CLK _17001_/D vssd1 vssd1 vccd1 vccd1 _17001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14213_ hold1505/X _14198_/B _14212_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ hold4966/X _12308_/B _11424_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11425_/X
+ sky130_fd_sc_hd__o211a_1
X_15193_ _15193_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ _15543_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14144_/Y sky130_fd_sc_hd__nand2_1
X_11356_ hold5250/X _11738_/B _11355_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ hold1941/X hold4925/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14075_ hold2467/X _14107_/A2 _14074_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14075_/X
+ sky130_fd_sc_hd__o211a_1
X_11287_ hold5623/X _11789_/B _11286_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13026_ hold990/X hold957/A _13043_/C vssd1 vssd1 vccd1 vccd1 _13028_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16312_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17903_ _17903_/CLK _17903_/D vssd1 vssd1 vccd1 vccd1 _17903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10238_ hold1513/X hold3789/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10239_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17479_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10169_ hold1757/X hold4617/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__mux2_1
X_17834_ _17834_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ hold5979/X _15004_/B hold938/X _15482_/A vssd1 vssd1 vccd1 vccd1 hold939/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17765_ _18003_/CLK _17765_/D vssd1 vssd1 vccd1 vccd1 _17765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _18305_/CLK _16716_/D vssd1 vssd1 vccd1 vccd1 _16716_/Q sky130_fd_sc_hd__dfxtp_1
X_13928_ hold246/X _17770_/Q hold124/X vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__mux2_1
XFILLER_0_187_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ _17696_/CLK _17696_/D vssd1 vssd1 vccd1 vccd1 _17696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _18205_/CLK _16647_/D vssd1 vssd1 vccd1 vccd1 _16647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13859_ _17740_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__and3_1
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16578_ _18166_/CLK _16578_/D vssd1 vssd1 vccd1 vccd1 _16578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18317_ _18349_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
X_15529_ _15529_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09050_ hold222/X hold489/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__mux2_1
X_18248_ _18376_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08001_ _14116_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__or2_1
X_18179_ _18199_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold513 hold513/A vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold524 input64/X vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__buf_1
XFILLER_0_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold535 hold535/A vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 hold546/A vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 hold557/A vssd1 vssd1 vccd1 vccd1 input50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 hold83/X vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__buf_4
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ hold4821/X _10049_/B _09951_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09952_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _12426_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _16069_/D sky130_fd_sc_hd__and2_1
XFILLER_0_216_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09883_ hold4733/X _10601_/B _09882_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09883_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _14438_/X vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ hold346/X hold434/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__mux2_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _15216_/X vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _08398_/X vssd1 vssd1 vccd1 vccd1 _15829_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 _16312_/Q vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _08396_/X vssd1 vssd1 vccd1 vccd1 _15828_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1257 _07889_/X vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ hold379/X hold775/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1268 _14418_/X vssd1 vssd1 vccd1 vccd1 _18005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1279 _18228_/Q vssd1 vssd1 vccd1 vccd1 hold1279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _12416_/A hold375/X vssd1 vssd1 vccd1 vccd1 _15969_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_400_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17887_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09317_ _15105_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09248_ _12759_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _16235_/D sky130_fd_sc_hd__and2_1
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09179_ hold733/X hold533/A vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__or2_2
XFILLER_0_44_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11210_ _11210_/A _11210_/B _11762_/C vssd1 vssd1 vccd1 vccd1 _11210_/X sky130_fd_sc_hd__and3_1
X_12190_ hold4946/X _12317_/B _12189_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _12190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11141_ _16871_/Q _11147_/B _11147_/C vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__and3_1
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput77 _13169_/A vssd1 vssd1 vccd1 vccd1 output77/X sky130_fd_sc_hd__buf_6
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ hold1644/X _16848_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__mux2_1
Xoutput88 _13249_/A vssd1 vssd1 vccd1 vccd1 output88/X sky130_fd_sc_hd__buf_6
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 _13097_/A vssd1 vssd1 vccd1 vccd1 output99/X sky130_fd_sc_hd__buf_6
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3160 _12581_/X vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _15185_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__or2_1
X_10023_ _13174_/A _11106_/A _10022_/X vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__a21oi_1
Xhold3171 _17499_/Q vssd1 vssd1 vccd1 vccd1 hold3171/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _17254_/CLK _15880_/D vssd1 vssd1 vccd1 vccd1 _15880_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3182 _12815_/X vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3193 _18329_/Q vssd1 vssd1 vccd1 vccd1 hold3193/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2470 _08253_/X vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ hold1170/X _14826_/B _14830_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14831_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2481 _14911_/X vssd1 vssd1 vccd1 vccd1 _18241_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 _18150_/Q vssd1 vssd1 vccd1 vccd1 hold2492/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _18215_/CLK _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1780 _09314_/X vssd1 vssd1 vccd1 vccd1 _16267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1791 _18216_/Q vssd1 vssd1 vccd1 vccd1 hold1791/X sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ _15209_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14762_/X sky130_fd_sc_hd__or2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ hold5465/X _13862_/B _11973_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11974_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _18350_/CLK _16501_/D vssd1 vssd1 vccd1 vccd1 _16501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13713_/A _13713_/B vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__or2_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ hold2681/X hold3810/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17481_ _17481_/CLK _17481_/D vssd1 vssd1 vccd1 vccd1 _17481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14693_ hold2850/X _14720_/B _14692_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16432_ _18377_/CLK _16432_/D vssd1 vssd1 vccd1 vccd1 _16432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_141_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18370_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13644_ _13761_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__or2_1
X_10856_ hold1042/X _16776_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16363_ _18346_/CLK _16363_/D vssd1 vssd1 vccd1 vccd1 _16363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13698_/A _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__or2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10787_ hold1534/X _16753_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _10788_/B sky130_fd_sc_hd__mux2_1
X_18102_ _18186_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15314_ _15344_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ hold2203/X hold3157/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__mux2_1
X_16294_ _16312_/CLK _16294_/D vssd1 vssd1 vccd1 vccd1 _16294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18033_ _18036_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
X_15245_ hold198/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12457_ hold17/X _12509_/A2 _12507_/A3 _12456_/X _09015_/A vssd1 vssd1 vccd1 vccd1
+ hold18/A sky130_fd_sc_hd__o311a_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ hold1420/X hold4399/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__mux2_1
X_15176_ hold2766/X _15167_/B _15175_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12388_ _15364_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _17287_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ hold2795/X _14148_/B _14126_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__o211a_1
X_11339_ hold2337/X _16937_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ hold915/X _14104_/B vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _14972_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17817_ _18425_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ hold163/X hold706/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold707/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_229_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17748_ _17748_/CLK _17748_/D vssd1 vssd1 vccd1 vccd1 _17748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08481_ hold1595/X _08486_/B _08480_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08481_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17679_ _17712_/CLK _17679_/D vssd1 vssd1 vccd1 vccd1 _17679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _15543_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09033_ _12430_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _16133_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 input16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold332 hold332/A vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__clkbuf_2
Xhold343 hold343/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold365/A vssd1 vssd1 vccd1 vccd1 input47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold376/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold387 hold387/A vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _15068_/A vssd1 vssd1 vccd1 vccd1 _15226_/C1 sky130_fd_sc_hd__buf_4
X_09935_ hold1983/X _16469_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__mux2_1
Xfanout812 _15026_/A vssd1 vssd1 vccd1 vccd1 _15192_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout823 _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__buf_4
XFILLER_0_217_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout834 fanout847/X vssd1 vssd1 vccd1 vccd1 _14805_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout845 _14815_/C1 vssd1 vssd1 vccd1 vccd1 _14865_/C1 sky130_fd_sc_hd__buf_4
Xfanout856 _15219_/A vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__buf_12
XFILLER_0_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09866_ _18357_/Q _16446_/Q _10034_/C vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__mux2_1
Xfanout867 _11203_/A vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__buf_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _08409_/X vssd1 vssd1 vccd1 vccd1 hold1010/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 _15199_/A vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__buf_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 _15043_/X vssd1 vssd1 vccd1 vccd1 _15044_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _14854_/A vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__buf_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _15142_/X vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ _09055_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1043 _18287_/Q vssd1 vssd1 vccd1 vccd1 hold1043/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _18378_/Q vssd1 vssd1 vccd1 vccd1 hold1054/X sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ hold2979/X hold3388/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__mux2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1065 hold1140/X vssd1 vssd1 vccd1 vccd1 hold1141/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 _18347_/Q vssd1 vssd1 vccd1 vccd1 hold1076/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _15414_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _15994_/D sky130_fd_sc_hd__and2_1
Xhold1087 _08426_/X vssd1 vssd1 vccd1 vccd1 _15843_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 _15666_/Q vssd1 vssd1 vccd1 vccd1 hold1098/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ hold596/X hold881/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold882/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10710_ _11121_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__or2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11690_ hold2197/X hold4469/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10641_ hold3571/X _10527_/A _10640_/X vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ hold4338/X _13856_/B _13359_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10572_ hold4616/X _10560_/A _10571_/X vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12311_ _17261_/Q _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ _13290_/X _16929_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15030_ _15030_/A _15030_/B vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__and2_1
X_12242_ hold2310/X _17238_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ hold2929/X hold4301/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11124_ _11124_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16981_ _18062_/CLK _16981_/D vssd1 vssd1 vccd1 vccd1 _16981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15932_ _17321_/CLK _15932_/D vssd1 vssd1 vccd1 vccd1 hold667/A sky130_fd_sc_hd__dfxtp_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11139_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10006_ _11158_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _16492_/D sky130_fd_sc_hd__nor2_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _17734_/CLK _15863_/D vssd1 vssd1 vccd1 vccd1 _15863_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_393_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17899_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14814_ _15099_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17666_/CLK _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _17722_/CLK _15794_/D vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_322_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17905_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ _18364_/CLK _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_1
X_14745_ hold2260/X _14772_/B _14744_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14745_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ hold1917/X hold4409/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10908_ _11115_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__or2_1
X_17464_ _17485_/CLK _17464_/D vssd1 vssd1 vccd1 vccd1 _17464_/Q sky130_fd_sc_hd__dfxtp_1
X_14676_ _15231_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14676_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ hold1353/X hold3320/X _13877_/C vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16415_ _18294_/CLK _16415_/D vssd1 vssd1 vccd1 vccd1 _16415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13627_ hold5709/X _13829_/B _13626_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13627_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17395_ _18445_/CLK _17395_/D vssd1 vssd1 vccd1 vccd1 _17395_/Q sky130_fd_sc_hd__dfxtp_1
X_10839_ _11694_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _18360_/CLK _16346_/D vssd1 vssd1 vccd1 vccd1 _16346_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ hold4135/X _13883_/B _13557_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ hold8/X _12509_/A2 _08868_/X _12508_/X _09015_/A vssd1 vssd1 vccd1 vccd1
+ hold9/A sky130_fd_sc_hd__o311a_1
XFILLER_0_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ _17510_/CLK _16277_/D vssd1 vssd1 vccd1 vccd1 _16277_/Q sky130_fd_sc_hd__dfxtp_1
X_13489_ hold4297/X _13777_/A2 _13488_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5309 _12139_/X vssd1 vssd1 vccd1 vccd1 _17203_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15228_ hold2691/X _15219_/B _15227_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15228_/X
+ sky130_fd_sc_hd__o211a_1
X_18016_ _18016_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4608 _16355_/Q vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4619 _16542_/Q vssd1 vssd1 vccd1 vccd1 hold4619/X sky130_fd_sc_hd__dlygate4sd3_1
X_15159_ _15213_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3907 _10477_/X vssd1 vssd1 vccd1 vccd1 _16649_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3918 _17189_/Q vssd1 vssd1 vccd1 vccd1 hold3918/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3929 _11242_/X vssd1 vssd1 vccd1 vccd1 _16904_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_205_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07981_ hold2256/X _07991_/A2 _07980_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09720_ _09936_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09651_ _09987_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08602_ _12426_/A hold894/X vssd1 vssd1 vccd1 vccd1 _15923_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09582_ _10482_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08533_ _12430_/A hold626/X vssd1 vssd1 vccd1 vccd1 _15890_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08464_ _14517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ _15509_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5810 output99/X vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_12
X_09016_ hold174/X hold543/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5821 output94/X vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_170_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5832 hold5832/A vssd1 vssd1 vccd1 vccd1 hold5832/X sky130_fd_sc_hd__buf_2
Xhold5843 _16282_/Q vssd1 vssd1 vccd1 vccd1 hold5843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5854 hold5854/A vssd1 vssd1 vccd1 vccd1 hold5854/X sky130_fd_sc_hd__buf_2
Xhold140 hold11/X vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__buf_4
Xhold5865 _16285_/Q vssd1 vssd1 vccd1 vccd1 hold5865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5876 hold5876/A vssd1 vssd1 vccd1 vccd1 hold5876/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold162 input36/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold173 input35/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5887 _18421_/Q vssd1 vssd1 vccd1 vccd1 hold5887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5898 _07826_/X vssd1 vssd1 vccd1 vccd1 hold5898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 _09349_/Y vssd1 vssd1 vccd1 vccd1 _15485_/A2 sky130_fd_sc_hd__buf_8
Xfanout631 _12445_/A vssd1 vssd1 vccd1 vccd1 _12509_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_217_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__or2_1
Xfanout642 _12807_/A vssd1 vssd1 vccd1 vccd1 _12789_/A sky130_fd_sc_hd__buf_2
Xfanout653 _12909_/A vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__clkbuf_4
Xfanout664 _12981_/A vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__buf_4
XFILLER_0_232_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout675 _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08369_/A sky130_fd_sc_hd__buf_4
Xfanout686 _14013_/C1 vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__buf_4
X_09849_ _11082_/A _09849_/B vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__or2_1
Xfanout697 _12396_/A vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12860_ hold3314/X _12859_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12861_/B sky130_fd_sc_hd__mux2_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11811_ _13797_/A _11811_/B vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__or2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12791_ hold3347/X _12790_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__mux2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ hold1634/X _14535_/B _14529_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14530_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ hold4681/X _12219_/A _11741_/X vssd1 vssd1 vccd1 vccd1 _11742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ _14910_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14461_/X sky130_fd_sc_hd__or2_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11694_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__or2_1
X_16200_ _17507_/CLK _16200_/D vssd1 vssd1 vccd1 vccd1 _16200_/Q sky130_fd_sc_hd__dfxtp_1
X_13412_ hold1245/X _17591_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__mux2_1
X_10624_ _11194_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _16698_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17180_ _17198_/CLK _17180_/D vssd1 vssd1 vccd1 vccd1 _17180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ _14392_/A _14392_/B vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16131_ _16131_/CLK _16131_/D vssd1 vssd1 vccd1 vccd1 hold429/A sky130_fd_sc_hd__dfxtp_1
X_13343_ hold2643/X hold5681/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__mux2_1
X_10555_ hold4923/X _10649_/B _10554_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16062_ _17297_/CLK _16062_/D vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _17585_/Q _17119_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__mux2_1
X_10486_ hold4721/X _10598_/B _10485_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ hold2654/X _15004_/B _15012_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15013_/X
+ sky130_fd_sc_hd__o211a_1
X_12225_ _13794_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12156_ _12231_/A _12156_/B vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ hold5593/X _11201_/B _11106_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _11107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12087_ _13461_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__or2_1
X_16964_ _17842_/CLK _16964_/D vssd1 vssd1 vccd1 vccd1 _16964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15915_ _18415_/CLK _15915_/D vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__dfxtp_1
X_11038_ hold4189/X _11729_/B _11037_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _11038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16895_ _18067_/CLK _16895_/D vssd1 vssd1 vccd1 vccd1 _16895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _17642_/CLK _15846_/D vssd1 vssd1 vccd1 vccd1 _15846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _17612_/CLK _15777_/D vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfxtp_1
X_12989_ hold3271/X _12988_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__mux2_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ _18398_/CLK _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14728_ _14782_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14659_ hold2953/X _14664_/B _14658_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14659_/X
+ sky130_fd_sc_hd__o211a_1
X_17447_ _17455_/CLK _17447_/D vssd1 vssd1 vccd1 vccd1 _17447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ hold2575/X _08209_/B _08179_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08180_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17378_ _17378_/CLK _17378_/D vssd1 vssd1 vccd1 vccd1 _17378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16329_ _18418_/CLK _16329_/D vssd1 vssd1 vccd1 vccd1 _16329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_24_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_24_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5106 _16902_/Q vssd1 vssd1 vccd1 vccd1 hold5106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5117 _11845_/X vssd1 vssd1 vccd1 vccd1 _17105_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5128 _17200_/Q vssd1 vssd1 vccd1 vccd1 hold5128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5139 _13339_/X vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4405 _17749_/Q vssd1 vssd1 vccd1 vccd1 hold4405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4416 _11050_/X vssd1 vssd1 vccd1 vccd1 _16840_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4427 _16860_/Q vssd1 vssd1 vccd1 vccd1 hold4427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4438 _11602_/X vssd1 vssd1 vccd1 vccd1 _17024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3704 _17720_/Q vssd1 vssd1 vccd1 vccd1 hold3704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4449 _17616_/Q vssd1 vssd1 vccd1 vccd1 hold4449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3715 _10498_/X vssd1 vssd1 vccd1 vccd1 _16656_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3726 _16607_/Q vssd1 vssd1 vccd1 vccd1 hold3726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3737 _12372_/Y vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3748 _16560_/Q vssd1 vssd1 vccd1 vccd1 hold3748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3759 _11148_/Y vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_244_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18210_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07964_ _15533_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09703_ hold3388/X _10025_/B _09702_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09703_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07895_ hold2162/X _07918_/B _07894_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _07895_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09634_ hold4481/X _09832_/A2 _09633_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _09634_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09565_ hold3631/X _10055_/B _09564_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08516_ hold1188/X _08503_/Y _08515_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ _09496_/A _15229_/A _15173_/A vssd1 vssd1 vccd1 vccd1 _09498_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_4_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_63_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_63_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ hold689/A hold732/A hold764/A hold752/A vssd1 vssd1 vccd1 vccd1 _14913_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08378_ hold367/X hold663/X hold134/X vssd1 vssd1 vccd1 vccd1 hold664/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ hold3130/X hold3718/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5640 _11860_/X vssd1 vssd1 vccd1 vccd1 _17110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ hold2689/X hold4897/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__mux2_1
Xhold5651 _11569_/X vssd1 vssd1 vccd1 vccd1 _17013_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5662 _09574_/X vssd1 vssd1 vccd1 vccd1 _16348_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5673 _16504_/Q vssd1 vssd1 vccd1 vccd1 hold5673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5684 _09688_/X vssd1 vssd1 vccd1 vccd1 _16386_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ hold4915/X _13811_/B _12009_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _12010_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4950 _16701_/Q vssd1 vssd1 vccd1 vccd1 hold4950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5695 _17602_/Q vssd1 vssd1 vccd1 vccd1 hold5695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4961 _11202_/Y vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4972 _17160_/Q vssd1 vssd1 vccd1 vccd1 hold4972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4983 _11587_/X vssd1 vssd1 vccd1 vccd1 _17019_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4994 _17255_/Q vssd1 vssd1 vccd1 vccd1 hold4994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout450 _11747_/C vssd1 vssd1 vccd1 vccd1 _12317_/C sky130_fd_sc_hd__clkbuf_8
Xfanout461 _12251_/S vssd1 vssd1 vccd1 vccd1 _12362_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 _11480_/S vssd1 vssd1 vccd1 vccd1 _11594_/S sky130_fd_sc_hd__buf_4
X_13961_ hold2331/X _13995_/A2 _13960_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _13961_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout483 _11147_/C vssd1 vssd1 vccd1 vccd1 _11156_/C sky130_fd_sc_hd__clkbuf_8
Xfanout494 _10025_/C vssd1 vssd1 vccd1 vccd1 _10001_/C sky130_fd_sc_hd__buf_6
XFILLER_0_214_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _17711_/CLK _15700_/D vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfxtp_1
X_12912_ _12912_/A _12912_/B vssd1 vssd1 vccd1 vccd1 _17480_/D sky130_fd_sc_hd__and2_1
X_16680_ _18144_/CLK _16680_/D vssd1 vssd1 vccd1 vccd1 _16680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ hold391/A hold532/X vssd1 vssd1 vccd1 vccd1 _14163_/B sky130_fd_sc_hd__or2_4
XFILLER_0_241_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _18428_/CLK _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
X_12843_ _12870_/A _12843_/B vssd1 vssd1 vccd1 vccd1 _17457_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18350_ _18350_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
X_15562_ _17898_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12780_/A _12774_/B vssd1 vssd1 vccd1 vccd1 _17434_/D sky130_fd_sc_hd__and2_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/CLK _17301_/D vssd1 vssd1 vccd1 vccd1 hold492/A sky130_fd_sc_hd__dfxtp_1
X_14513_ _15193_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__or2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ _12310_/A _11725_/B vssd1 vssd1 vccd1 vccd1 _17065_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18281_ _18351_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
X_15493_ _15509_/A _18424_/Q hold691/X vssd1 vssd1 vccd1 vccd1 _15493_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14444_ hold1406/X _14433_/B _14443_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14444_/X
+ sky130_fd_sc_hd__o211a_1
X_17232_ _17718_/CLK _17232_/D vssd1 vssd1 vccd1 vccd1 _17232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11656_ hold5605/X _11753_/B _11655_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _16693_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__and3_1
X_17163_ _17195_/CLK _17163_/D vssd1 vssd1 vccd1 vccd1 _17163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14375_ hold246/X _17985_/Q hold333/X vssd1 vssd1 vccd1 vccd1 hold334/A sky130_fd_sc_hd__mux2_1
XFILLER_0_141_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ hold4982/X _12317_/B _11586_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _17339_/CLK _16114_/D vssd1 vssd1 vccd1 vccd1 hold516/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _13800_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__or2_1
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ hold2180/X _16670_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__mux2_1
X_17094_ _17719_/CLK _17094_/D vssd1 vssd1 vccd1 vccd1 _17094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16045_ _17301_/CLK _16045_/D vssd1 vssd1 vccd1 vccd1 hold615/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13257_ _13257_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__and2_1
X_10469_ hold1170/X _16647_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12208_ hold5006/X _13811_/B _12207_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__o211a_1
X_13188_ hold4614/X _13187_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ hold5308/X _12329_/B _12138_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _12139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17996_ _17996_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1609 _15704_/Q vssd1 vssd1 vccd1 vccd1 hold1609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16947_ _17825_/CLK _16947_/D vssd1 vssd1 vccd1 vccd1 _16947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16878_ _18337_/CLK _16878_/D vssd1 vssd1 vccd1 vccd1 _16878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15829_ _17725_/CLK _15829_/D vssd1 vssd1 vccd1 vccd1 _15829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _15543_/A _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09360_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_75_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08301_ _15199_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _15557_/A hold1686/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08232_ hold915/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08163_ _08163_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _15719_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08094_ _15553_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4202 _12031_/X vssd1 vssd1 vccd1 vccd1 _17167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4213 _17690_/Q vssd1 vssd1 vccd1 vccd1 hold4213/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_425_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17179_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4224 _10852_/X vssd1 vssd1 vccd1 vccd1 _16774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4235 _17204_/Q vssd1 vssd1 vccd1 vccd1 hold4235/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3501 _13780_/X vssd1 vssd1 vccd1 vccd1 _17713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4246 _13789_/X vssd1 vssd1 vccd1 vccd1 _17716_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3512 _13678_/X vssd1 vssd1 vccd1 vccd1 _17679_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4257 _17214_/Q vssd1 vssd1 vccd1 vccd1 hold4257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4268 _12172_/X vssd1 vssd1 vccd1 vccd1 _17214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3523 _16991_/Q vssd1 vssd1 vccd1 vccd1 hold3523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3534 _11059_/X vssd1 vssd1 vccd1 vccd1 _16843_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4279 _16774_/Q vssd1 vssd1 vccd1 vccd1 hold4279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3545 _16530_/Q vssd1 vssd1 vccd1 vccd1 hold3545/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2800 _15653_/Q vssd1 vssd1 vccd1 vccd1 hold2800/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2811 _14542_/X vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3556 _10623_/Y vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08996_ _09015_/A hold499/X vssd1 vssd1 vccd1 vccd1 _16115_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3567 _16912_/Q vssd1 vssd1 vccd1 vccd1 hold3567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2822 _14031_/X vssd1 vssd1 vccd1 vccd1 _17819_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3578 _12608_/X vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 _09173_/X vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2844 _18445_/Q vssd1 vssd1 vccd1 vccd1 hold2844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3589 hold4052/X vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 _14023_/X vssd1 vssd1 vccd1 vccd1 _17815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2866 _14787_/X vssd1 vssd1 vccd1 vccd1 _18182_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07947_ hold2645/X _07978_/B _07946_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2877 _09334_/X vssd1 vssd1 vccd1 vccd1 _16277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2888 _17781_/Q vssd1 vssd1 vccd1 vccd1 hold2888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2899 _17967_/Q vssd1 vssd1 vccd1 vccd1 hold2899/X sky130_fd_sc_hd__dlygate4sd3_1
X_07878_ hold2658/X _07865_/B _07877_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _07878_/X
+ sky130_fd_sc_hd__o211a_1
X_09617_ _18274_/Q hold3422/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ hold3168/X _13190_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09479_ hold850/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09481_/C sky130_fd_sc_hd__or2_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ hold2467/X _16994_/Q _12344_/C vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ _17338_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ hold2939/X hold4103/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ hold808/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__or2_1
X_11372_ hold2925/X _16948_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11373_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13111_ _13199_/A1 _13109_/X _13110_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13111_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_46_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10323_ _10497_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14091_ hold2068/X _14094_/B _14090_/Y _12975_/A vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_166_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _13046_/C _13046_/D hold932/X vssd1 vssd1 vccd1 vccd1 hold933/A sky130_fd_sc_hd__nor3_1
Xhold5470 _11689_/X vssd1 vssd1 vccd1 vccd1 _17053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10254_ _10536_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__or2_1
Xhold5481 _16773_/Q vssd1 vssd1 vccd1 vccd1 hold5481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5492 _10870_/X vssd1 vssd1 vccd1 vccd1 _16780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4780 _12357_/Y vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17850_ _18425_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10185_ _10560_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__or2_1
Xhold4791 _16556_/Q vssd1 vssd1 vccd1 vccd1 hold4791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16801_ _18068_/CLK _16801_/D vssd1 vssd1 vccd1 vccd1 _16801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17781_ _17816_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_1
X_14993_ hold2995/X hold514/X _14992_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _14993_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout280 _12273_/A vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__buf_4
Xfanout291 _12051_/A vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__buf_2
XFILLER_0_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16732_ _17997_/CLK _16732_/D vssd1 vssd1 vccd1 vccd1 _16732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13944_ _15559_/A hold1525/X hold124/X vssd1 vssd1 vccd1 vccd1 _13944_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16663_ _18123_/CLK _16663_/D vssd1 vssd1 vccd1 vccd1 _16663_/Q sky130_fd_sc_hd__dfxtp_1
X_13875_ hold3312/X _13788_/A _13874_/X vssd1 vssd1 vccd1 vccd1 _13875_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18402_ _18402_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
X_15614_ _17113_/CLK _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_12826_ hold2347/X _17453_/Q _12826_/S vssd1 vssd1 vccd1 vccd1 _12826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16594_ _18208_/CLK _16594_/D vssd1 vssd1 vccd1 vccd1 _16594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ _18389_/CLK hold384/X vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
X_12757_ hold2784/X _17430_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__mux2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15545_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ hold2594/X _17060_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__mux2_1
X_18264_ _18296_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
X_15476_ hold397/X _09392_/B _09386_/D hold438/X _15475_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_189_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12688_ hold1947/X _17407_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14427_ _15541_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17215_ _17215_/CLK _17215_/D vssd1 vssd1 vccd1 vccd1 _17215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11639_ hold1472/X _17037_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__mux2_1
X_18195_ _18227_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ _14360_/A _14358_/B vssd1 vssd1 vccd1 vccd1 _17976_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17146_ _17178_/CLK _17146_/D vssd1 vssd1 vccd1 vccd1 _17146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold706 hold706/A vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 input53/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 hold728/A vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _13308_/X hold4617/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17077_ _17901_/CLK _17077_/D vssd1 vssd1 vccd1 vccd1 _17077_/Q sky130_fd_sc_hd__dfxtp_1
Xhold739 hold739/A vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ hold1958/X hold756/X _14288_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14289_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ _17284_/CLK _16028_/D vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08850_ hold263/X hold737/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold738/A sky130_fd_sc_hd__mux2_1
Xhold2107 _15682_/Q vssd1 vssd1 vccd1 vccd1 hold2107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2118 _15697_/Q vssd1 vssd1 vccd1 vccd1 hold2118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2129 _08430_/X vssd1 vssd1 vccd1 vccd1 _15845_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07801_ _09342_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__and2_1
Xhold1406 _18018_/Q vssd1 vssd1 vccd1 vccd1 hold1406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08781_ hold222/X hold385/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold386/A sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1417 _14506_/X vssd1 vssd1 vccd1 vccd1 _18047_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _18430_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1428 _07901_/X vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 hold1439/A vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09402_ _12404_/A _09402_/B vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__and2_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _15555_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09264_ _12738_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _16243_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _15549_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08215_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09195_ hold1166/X _09218_/B _09194_/X _12807_/A vssd1 vssd1 vccd1 vccd1 _09195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _14330_/A hold1353/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ hold1363/X _08097_/A2 _08076_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _08077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4010 _17626_/Q vssd1 vssd1 vccd1 vccd1 hold4010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4021 _09604_/X vssd1 vssd1 vccd1 vccd1 _16358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4032 _17627_/Q vssd1 vssd1 vccd1 vccd1 hold4032/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4043 _10168_/X vssd1 vssd1 vccd1 vccd1 _16546_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4054 _10420_/X vssd1 vssd1 vccd1 vccd1 _16630_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3320 _17120_/Q vssd1 vssd1 vccd1 vccd1 hold3320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4065 _16642_/Q vssd1 vssd1 vccd1 vccd1 hold4065/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4076 _10552_/X vssd1 vssd1 vccd1 vccd1 _16674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3331 _17389_/Q vssd1 vssd1 vccd1 vccd1 hold3331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4087 _17140_/Q vssd1 vssd1 vccd1 vccd1 hold4087/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3342 _17437_/Q vssd1 vssd1 vccd1 vccd1 hold3342/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4098 _09694_/X vssd1 vssd1 vccd1 vccd1 _16388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3353 _17453_/Q vssd1 vssd1 vccd1 vccd1 hold3353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3364 _09898_/X vssd1 vssd1 vccd1 vccd1 _16456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__buf_4
XFILLER_0_216_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3375 _16489_/Q vssd1 vssd1 vccd1 vccd1 hold3375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2630 _16167_/Q vssd1 vssd1 vccd1 vccd1 hold2630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3386 _16435_/Q vssd1 vssd1 vccd1 vccd1 hold3386/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2641 _07969_/X vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ hold607/X hold656/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold657/A sky130_fd_sc_hd__mux2_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_4
Xhold2652 _18109_/Q vssd1 vssd1 vccd1 vccd1 hold2652/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3397 _17457_/Q vssd1 vssd1 vccd1 vccd1 hold3397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2663 _16242_/Q vssd1 vssd1 vccd1 vccd1 hold2663/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2674 _15765_/Q vssd1 vssd1 vccd1 vccd1 hold2674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 _18264_/Q vssd1 vssd1 vccd1 vccd1 hold2685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1940 _14219_/X vssd1 vssd1 vccd1 vccd1 _17909_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__buf_4
Xhold1951 _14611_/X vssd1 vssd1 vccd1 vccd1 _18097_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__buf_4
Xhold2696 _15230_/X vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ hold2459/X hold4085/X _13556_/S vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__mux2_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1962 _18159_/Q vssd1 vssd1 vccd1 vccd1 hold1962/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1973 _17891_/Q vssd1 vssd1 vccd1 vccd1 hold1973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 _15200_/X vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1995 _14931_/X vssd1 vssd1 vccd1 vccd1 _18250_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _11637_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13660_ hold4391/X _13880_/B _13659_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13660_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _11064_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ hold3610/X _12610_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ hold3458/X _13880_/B _13590_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13591_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15330_ hold335/X _15486_/A2 _09357_/B hold314/X vssd1 vssd1 vccd1 vccd1 _15330_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ hold3257/X _12541_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15261_ _16290_/Q _15477_/A2 _15487_/B1 _16078_/Q _15260_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12473_ hold74/X _12445_/A _12445_/B _12472_/X _12436_/A vssd1 vssd1 vccd1 vccd1
+ hold75/A sky130_fd_sc_hd__o311a_1
XFILLER_0_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_347_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17737_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17000_ _18427_/CLK _17000_/D vssd1 vssd1 vccd1 vccd1 _17000_/Q sky130_fd_sc_hd__dfxtp_1
X_14212_ _15557_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or2_1
X_11424_ _12213_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ hold2250/X _15219_/B _15191_/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 _15192_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_8 _13156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14143_ hold2508/X _14142_/B _14142_/Y _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14143_/X
+ sky130_fd_sc_hd__o211a_1
X_11355_ _11643_/A _11355_/B vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ hold3764/X _10628_/B _10305_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10306_/X
+ sky130_fd_sc_hd__o211a_1
X_14074_ _14862_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14074_/X sky130_fd_sc_hd__or2_1
X_11286_ _11670_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13025_ hold958/X _13025_/B _13025_/C vssd1 vssd1 vccd1 vccd1 _17518_/D sky130_fd_sc_hd__and3_1
X_17902_ _17902_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10237_ hold5381/X _10619_/B _10236_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17833_ _17842_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_1
X_10168_ hold4042/X _10622_/B _10167_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10168_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17764_ _17935_/CLK _17764_/D vssd1 vssd1 vccd1 vccd1 _17764_/Q sky130_fd_sc_hd__dfxtp_1
X_10099_ hold3689/X _10601_/B _10098_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14976_ hold926/X _15018_/B vssd1 vssd1 vccd1 vccd1 hold938/A sky130_fd_sc_hd__or2_1
XFILLER_0_234_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16715_ _18045_/CLK _16715_/D vssd1 vssd1 vccd1 vccd1 _16715_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_63_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18006_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13927_ _13927_/A hold698/X vssd1 vssd1 vccd1 vccd1 _17769_/D sky130_fd_sc_hd__and2_1
X_17695_ _17695_/CLK _17695_/D vssd1 vssd1 vccd1 vccd1 _17695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646_ _18202_/CLK _16646_/D vssd1 vssd1 vccd1 vccd1 _16646_/Q sky130_fd_sc_hd__dfxtp_1
X_13858_ _13873_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _17739_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ hold3330/X _12808_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_169_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16577_ _18229_/CLK _16577_/D vssd1 vssd1 vccd1 vccd1 _16577_/Q sky130_fd_sc_hd__dfxtp_1
X_13789_ hold4245/X _13883_/B _13788_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18316_ _18316_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ hold1125/X _15547_/B _15527_/X _12759_/A vssd1 vssd1 vccd1 vccd1 _15528_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _18389_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
X_15459_ hold265/X _09386_/A _09357_/A _17321_/Q _15458_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_167_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ hold1761/X _08033_/B _07999_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _08000_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18178_ _18178_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 hold503/A vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__buf_6
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17129_ _17129_/CLK _17129_/D vssd1 vssd1 vccd1 vccd1 _17129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold525 hold525/A vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__buf_8
XFILLER_0_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold536 hold536/A vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold547 hold547/A vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09951_ _09954_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__or2_1
Xhold558 input50/X vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__clkbuf_2
Xhold569 hold569/A vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ hold256/X hold442/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09882_ _10488_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__or2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08833_ _15344_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _16035_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _16235_/Q vssd1 vssd1 vccd1 vccd1 hold1203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 _18232_/Q vssd1 vssd1 vccd1 vccd1 hold1214/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1225 _15833_/Q vssd1 vssd1 vccd1 vccd1 hold1225/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1236 _09417_/X vssd1 vssd1 vccd1 vccd1 _16294_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _15374_/A hold257/X vssd1 vssd1 vccd1 vccd1 _16002_/D sky130_fd_sc_hd__and2_1
Xhold1247 hold1275/X vssd1 vssd1 vccd1 vccd1 hold1276/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1258 _15660_/Q vssd1 vssd1 vccd1 vccd1 hold1258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1269 _15587_/Q vssd1 vssd1 vccd1 vccd1 hold1269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ hold346/X hold374/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold375/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ hold3045/X _09325_/B _09315_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _15523_/A hold1203/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_440_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ hold733/X hold533/X vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08145_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _15703_/D sky130_fd_sc_hd__and2_1
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ hold3438/X _11729_/B _11139_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _11140_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 _13177_/A vssd1 vssd1 vccd1 vccd1 output78/X sky130_fd_sc_hd__buf_6
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ hold3974/X _11168_/B _11070_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _11071_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 _13257_/A vssd1 vssd1 vccd1 vccd1 output89/X sky130_fd_sc_hd__buf_6
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3150 _12875_/X vssd1 vssd1 vccd1 vccd1 _12876_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10022_ _16498_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__and3_1
Xhold3161 _17478_/Q vssd1 vssd1 vccd1 vccd1 hold3161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3172 _12968_/X vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3183 _17447_/Q vssd1 vssd1 vccd1 vccd1 hold3183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3194 _15094_/X vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2460 _08002_/X vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ hold972/X _14830_/B vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__or2_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2471 _15679_/Q vssd1 vssd1 vccd1 vccd1 hold2471/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 _15850_/Q vssd1 vssd1 vccd1 vccd1 hold2482/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 _14721_/X vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 _14229_/X vssd1 vssd1 vccd1 vccd1 _17914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ hold3084/X _14772_/B _14760_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14761_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1781 _18046_/Q vssd1 vssd1 vccd1 vccd1 hold1781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11973_ _12261_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__or2_1
Xhold1792 _14859_/X vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _18321_/CLK _16500_/D vssd1 vssd1 vccd1 vccd1 _16500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ hold2650/X hold3428/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13713_/B sky130_fd_sc_hd__mux2_1
X_10924_ hold4380/X _11210_/B _10923_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _10924_/X
+ sky130_fd_sc_hd__o211a_1
X_14692_ _15193_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__or2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17481_/CLK _17480_/D vssd1 vssd1 vccd1 vccd1 _17480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16431_ _18342_/CLK _16431_/D vssd1 vssd1 vccd1 vccd1 _16431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10855_ hold4283/X _11147_/B _10854_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10855_/X
+ sky130_fd_sc_hd__o211a_1
X_13643_ hold1755/X hold4559/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16362_ _18273_/CLK _16362_/D vssd1 vssd1 vccd1 vccd1 _16362_/Q sky130_fd_sc_hd__dfxtp_1
X_13574_ hold2723/X hold5282/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13575_/B sky130_fd_sc_hd__mux2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ hold4215/X _11732_/B _10785_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10786_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18101_ _18230_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15481_/A1 _15305_/X _15312_/X _15490_/B1 hold4585/X vssd1 vssd1 vccd1 vccd1
+ _15313_/X sky130_fd_sc_hd__a32o_1
X_12525_ _12531_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _17351_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16293_ _16311_/CLK _16293_/D vssd1 vssd1 vccd1 vccd1 _16293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_181_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18293_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032_ _18032_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
X_12456_ _17321_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__or2_1
X_15244_ _15264_/A _15244_/B vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__and2_1
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_110_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17332_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ hold3523/X _12344_/B _11406_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11407_/X
+ sky130_fd_sc_hd__o211a_1
X_15175_ _15229_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or2_1
X_12387_ hold113/X hold629/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _15525_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__or2_1
X_11338_ hold3932/X _12299_/B _11337_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ hold1561/X _14107_/A2 _14056_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14057_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11269_ hold5208/X _12314_/B _11268_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ hold1179/X _13003_/Y _13007_/X _15264_/A vssd1 vssd1 vccd1 vccd1 _13008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ _17816_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17747_ _17747_/CLK _17747_/D vssd1 vssd1 vccd1 vccd1 _17747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14959_ hold2685/X _14946_/B _14958_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08480_ _15213_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08480_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ _17680_/CLK _17678_/D vssd1 vssd1 vccd1 vccd1 _17678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16629_ _18193_/CLK _16629_/D vssd1 vssd1 vccd1 vccd1 _16629_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_269_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18182_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ hold2393/X _09106_/B _09100_/Y _12975_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09032_ hold256/X hold288/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 input16/X vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__buf_12
Xhold344 hold40/X vssd1 vssd1 vccd1 vccd1 input11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 input47/X vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold377 hold52/X vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold388 la_data_in[31] vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _10028_/A _10010_/B _09933_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09934_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout813 _15062_/A vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__buf_4
Xfanout824 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14879_/C1 sky130_fd_sc_hd__buf_4
Xfanout835 _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14835_/C1 sky130_fd_sc_hd__buf_4
Xfanout846 fanout847/X vssd1 vssd1 vccd1 vccd1 _14815_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09865_ hold4749/X _10055_/B _09864_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09865_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout857 _15221_/A vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__buf_12
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 _08160_/X vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 fanout873/X vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__clkbuf_16
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout879 _15199_/A vssd1 vssd1 vccd1 vccd1 hold1725/A sky130_fd_sc_hd__buf_6
Xhold1011 _08410_/X vssd1 vssd1 vccd1 vccd1 _15835_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _15044_/X vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ hold47/X hold701/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__mux2_1
Xhold1033 la_data_in[6] vssd1 vssd1 vccd1 vccd1 hold1033/X sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ hold5040/X _10034_/B _09795_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09796_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1044 _15007_/X vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _15196_/X vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1066 hold1142/X vssd1 vssd1 vccd1 vccd1 hold1066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _15132_/X vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ hold174/X hold198/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__mux2_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 _15881_/Q vssd1 vssd1 vccd1 vccd1 hold1088/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _08053_/X vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _09053_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _15960_/D sky130_fd_sc_hd__and2_1
XFILLER_0_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _16704_/Q _10646_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10571_ _10571_/A _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _17260_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13290_ _17587_/Q _17121_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ _12335_/A _12274_/A2 _12240_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12172_ hold4267/X _13871_/B _12171_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12172_/X
+ sky130_fd_sc_hd__o211a_1
X_11123_ hold2349/X hold4531/X _11219_/C vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16980_ _17858_/CLK _16980_/D vssd1 vssd1 vccd1 vccd1 _16980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15931_ _17347_/CLK _15931_/D vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__dfxtp_1
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ hold2814/X _16842_/Q _11150_/C vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__mux2_1
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ _13126_/A _09987_/A _10004_/X vssd1 vssd1 vccd1 vccd1 _10005_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _17739_/CLK _15862_/D vssd1 vssd1 vccd1 vccd1 _15862_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2290 _15813_/Q vssd1 vssd1 vccd1 vccd1 hold2290/X sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _17728_/CLK _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14813_ hold1094/X _14828_/B _14812_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _18447_/CLK _15793_/D vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17532_ _17534_/CLK _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14744_ _15191_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ hold5473/X _12052_/A2 _11955_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11956_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10907_ hold1837/X _16793_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__mux2_1
X_17463_ _17483_/CLK _17463_/D vssd1 vssd1 vccd1 vccd1 _17463_/Q sky130_fd_sc_hd__dfxtp_1
X_14675_ hold2341/X _14666_/B _14674_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14675_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_362_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17245_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ hold4519/X _12344_/B _11886_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__o211a_1
X_16414_ _18383_/CLK _16414_/D vssd1 vssd1 vccd1 vccd1 _16414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ _13734_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ hold3232/X hold5563/X _11768_/C vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__mux2_1
X_17394_ _18445_/CLK _17394_/D vssd1 vssd1 vccd1 vccd1 _17394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _18350_/CLK _16345_/D vssd1 vssd1 vccd1 vccd1 _16345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ hold2957/X _16747_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ _13788_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _17347_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__or2_1
Xclkbuf_6_14_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_14_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16276_ _17517_/CLK _16276_/D vssd1 vssd1 vccd1 vccd1 _16276_/Q sky130_fd_sc_hd__dfxtp_1
X_13488_ _13776_/A _13488_/B vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ _18016_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12439_ hold292/X hold598/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__mux2_1
X_15227_ _15227_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15227_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4609 _10074_/Y vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ hold1819/X _15165_/B _15157_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _15158_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3908 _16620_/Q vssd1 vssd1 vccd1 vccd1 hold3908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3919 _12001_/X vssd1 vssd1 vccd1 vccd1 _17157_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14109_ _14789_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14140_/B sky130_fd_sc_hd__or2_4
XFILLER_0_103_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15089_ _15197_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07980_ _15549_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ hold966/X _16374_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08601_ hold312/X hold893/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold894/A sky130_fd_sc_hd__mux2_1
XFILLER_0_207_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09581_ hold984/X _13278_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08532_ hold554/X hold625/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold626/A sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_53_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_53_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_08463_ hold2297/X _08488_/B _08462_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08463_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08394_ hold203/X hold754/X vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__or2_4
XFILLER_0_169_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09015_ _09015_/A hold597/X vssd1 vssd1 vccd1 vccd1 _16124_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5800 output81/X vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_12
Xhold5811 hold5945/X vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__buf_1
XFILLER_0_147_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5822 hold5949/X vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__buf_1
XFILLER_0_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5833 hold5965/X vssd1 vssd1 vccd1 vccd1 hold5833/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5844 hold5844/A vssd1 vssd1 vccd1 vccd1 hold5844/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold130 hold761/X vssd1 vssd1 vccd1 vccd1 hold762/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5855 _16283_/Q vssd1 vssd1 vccd1 vccd1 hold5855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5866 hold5866/A vssd1 vssd1 vccd1 vccd1 hold5866/X sky130_fd_sc_hd__clkbuf_4
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5877 hold6016/X vssd1 vssd1 vccd1 vccd1 hold5877/X sky130_fd_sc_hd__buf_2
Xhold163 hold65/X vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__buf_4
Xhold5888 hold5888/A vssd1 vssd1 vccd1 vccd1 hold5888/X sky130_fd_sc_hd__clkbuf_4
Xhold5899 hold6027/X vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__clkbuf_2
Xhold174 hold26/X vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__buf_4
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _09362_/C vssd1 vssd1 vccd1 vccd1 _15448_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_217_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout621 _09349_/Y vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__clkbuf_8
Xfanout632 _08597_/Y vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__clkbuf_8
X_09917_ hold856/X _16463_/Q _10019_/C vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout643 _12807_/A vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__buf_4
Xfanout654 _12909_/A vssd1 vssd1 vccd1 vccd1 _12912_/A sky130_fd_sc_hd__buf_4
Xfanout665 fanout693/X vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout676 fanout692/X vssd1 vssd1 vccd1 vccd1 _13672_/C1 sky130_fd_sc_hd__clkbuf_4
X_09848_ hold3029/X hold5038/X _11177_/C vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__mux2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 _14013_/C1 vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__buf_4
Xfanout698 _12386_/A vssd1 vssd1 vccd1 vccd1 _12531_/A sky130_fd_sc_hd__buf_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ hold1985/X _16417_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__mux2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ hold2506/X _17094_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ hold1166/X hold3177/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _17071_/Q _12314_/B _12314_/C vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__and3_1
XFILLER_0_230_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14460_ hold2721/X _14482_/A2 _14459_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14460_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ hold2514/X hold4360/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ hold3555/X _10527_/A _10622_/X vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__a21oi_1
X_13411_ hold5459/X _12353_/B _13410_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _13411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14391_ _15233_/A hold2647/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16130_ _18423_/CLK _16130_/D vssd1 vssd1 vccd1 vccd1 hold674/A sky130_fd_sc_hd__dfxtp_1
X_13342_ hold5689/X _13829_/B _13341_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__o211a_1
X_10554_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _13273_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13273_/X sky130_fd_sc_hd__and2_1
XFILLER_0_228_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ _18407_/CLK _16061_/D vssd1 vssd1 vccd1 vccd1 _16061_/Q sky130_fd_sc_hd__dfxtp_1
X_10485_ _10563_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _15227_/A _15016_/B vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__or2_1
X_12224_ hold2729/X hold5272/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ hold2201/X _17209_/Q _12251_/S vssd1 vssd1 vccd1 vccd1 _12156_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11106_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11106_/X sky130_fd_sc_hd__or2_1
X_12086_ hold2225/X _17186_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16963_ _17870_/CLK _16963_/D vssd1 vssd1 vccd1 vccd1 _16963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15914_ _17297_/CLK _15914_/D vssd1 vssd1 vccd1 vccd1 hold648/A sky130_fd_sc_hd__dfxtp_1
X_11037_ _11637_/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11037_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16894_ _17892_/CLK _16894_/D vssd1 vssd1 vccd1 vccd1 _16894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _17738_/CLK _15845_/D vssd1 vssd1 vccd1 vccd1 _15845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _17707_/CLK _15776_/D vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ hold1252/X _17507_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_235_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17515_ _17515_/CLK _17515_/D vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ hold2826/X _14714_/B _14726_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14727_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11939_ hold2824/X _17137_/Q _12314_/C vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17446_ _17446_/CLK _17446_/D vssd1 vssd1 vccd1 vccd1 _17446_/Q sky130_fd_sc_hd__dfxtp_1
X_14658_ _15105_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ hold3706/X _13814_/B _13608_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__o211a_1
X_17377_ _17517_/CLK _17377_/D vssd1 vssd1 vccd1 vccd1 _17377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ hold1956/X _14612_/B _14588_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14589_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16328_ _18413_/CLK _16328_/D vssd1 vssd1 vccd1 vccd1 _16328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5107 _11716_/X vssd1 vssd1 vccd1 vccd1 _17062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5118 _16486_/Q vssd1 vssd1 vccd1 vccd1 hold5118/X sky130_fd_sc_hd__dlygate4sd3_1
X_16259_ _17379_/CLK _16259_/D vssd1 vssd1 vccd1 vccd1 _16259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5129 _12034_/X vssd1 vssd1 vccd1 vccd1 _17168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4406 _13792_/X vssd1 vssd1 vccd1 vccd1 _17717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4417 _17239_/Q vssd1 vssd1 vccd1 vccd1 hold4417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4428 _11014_/X vssd1 vssd1 vccd1 vccd1 _16828_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4439 _16995_/Q vssd1 vssd1 vccd1 vccd1 hold4439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3705 _13705_/X vssd1 vssd1 vccd1 vccd1 _17688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3716 _16619_/Q vssd1 vssd1 vccd1 vccd1 hold3716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3727 _10255_/X vssd1 vssd1 vccd1 vccd1 _16575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3738 _17587_/Q vssd1 vssd1 vccd1 vccd1 hold3738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3749 _10114_/X vssd1 vssd1 vccd1 vccd1 _16528_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ hold2335/X _07978_/B _07962_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _07963_/X
+ sky130_fd_sc_hd__o211a_1
X_09702_ _09984_/A _09702_/B vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07894_ _14403_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09633_ _09843_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_284_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18052_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_213_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16517_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08515_ _15519_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__or2_1
X_09495_ _14555_/B _14555_/C _09495_/C vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__or3_1
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08446_ hold1487/X _08433_/B _08445_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _08377_/A hold206/X vssd1 vssd1 vccd1 vccd1 _15820_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5630 _11674_/X vssd1 vssd1 vccd1 vccd1 _17048_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10270_ hold3687/X _11180_/B _10269_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10270_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5641 _17077_/Q vssd1 vssd1 vccd1 vccd1 hold5641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5652 _16344_/Q vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5663 _17569_/Q vssd1 vssd1 vccd1 vccd1 hold5663/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5674 _09946_/X vssd1 vssd1 vccd1 vccd1 _16472_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5685 _17662_/Q vssd1 vssd1 vccd1 vccd1 hold5685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4940 _17226_/Q vssd1 vssd1 vccd1 vccd1 hold4940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4951 _10537_/X vssd1 vssd1 vccd1 vccd1 _16669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5696 _13351_/X vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4962 _16733_/Q vssd1 vssd1 vccd1 vccd1 hold4962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4973 _11914_/X vssd1 vssd1 vccd1 vccd1 _17128_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4984 _16915_/Q vssd1 vssd1 vccd1 vccd1 hold4984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4995 _12199_/X vssd1 vssd1 vccd1 vccd1 _17223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout440 _12029_/S vssd1 vssd1 vccd1 vccd1 _13817_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout451 _11747_/C vssd1 vssd1 vccd1 vccd1 _12314_/C sky130_fd_sc_hd__buf_6
XFILLER_0_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout462 _12251_/S vssd1 vssd1 vccd1 vccd1 _13868_/C sky130_fd_sc_hd__clkbuf_8
Xfanout473 _11204_/C vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__buf_6
X_13960_ _15521_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13960_/X sky130_fd_sc_hd__or2_1
Xfanout484 _11057_/S vssd1 vssd1 vccd1 vccd1 _11147_/C sky130_fd_sc_hd__buf_6
Xfanout495 _11096_/S vssd1 vssd1 vccd1 vccd1 _11192_/C sky130_fd_sc_hd__clkbuf_8
X_12911_ hold3390/X _12910_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ hold391/A hold532/X vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__nor2_1
XFILLER_0_216_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15630_ _17194_/CLK _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ hold3397/X _12841_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__mux2_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _17261_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ hold3778/X _12772_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17306_/CLK _17300_/D vssd1 vssd1 vccd1 vccd1 hold780/A sky130_fd_sc_hd__dfxtp_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ hold2147/X _14535_/B _14511_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14512_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18280_ _18374_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11724_ hold3579/X _11631_/A _11723_/X vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15492_ hold690/X hold122/X vssd1 vssd1 vccd1 vccd1 hold691/A sky130_fd_sc_hd__nand2_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17231_ _17263_/CLK _17231_/D vssd1 vssd1 vccd1 vccd1 _17231_/Q sky130_fd_sc_hd__dfxtp_1
X_14443_ _14443_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__or2_1
X_11655_ _11658_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10606_ _18461_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _16692_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_88_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18398_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17162_ _17194_/CLK _17162_/D vssd1 vssd1 vccd1 vccd1 _17162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11586_ _12285_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__or2_1
X_14374_ _14374_/A hold646/X vssd1 vssd1 vccd1 vccd1 _17984_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ _17340_/CLK _16113_/D vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10537_ hold4950/X _10631_/B _10536_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10537_/X
+ sky130_fd_sc_hd__o211a_1
X_13325_ hold2056/X hold3565/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17093_ _17253_/CLK _17093_/D vssd1 vssd1 vccd1 vccd1 _17093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16044_ _16128_/CLK _16044_/D vssd1 vssd1 vccd1 vccd1 hold737/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13256_ _13249_/X _13255_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_204_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10468_ hold4195/X _10468_/A2 _10467_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _10468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12288_/A _12207_/B vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13187_ _13186_/X _16916_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__mux2_1
X_10399_ hold3797/X _10649_/B _10398_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10399_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _12234_/A _12138_/B vssd1 vssd1 vccd1 vccd1 _12138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17995_ _18030_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12069_ _12261_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
X_16946_ _17884_/CLK _16946_/D vssd1 vssd1 vccd1 vccd1 _16946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16877_ _18016_/CLK _16877_/D vssd1 vssd1 vccd1 vccd1 _16877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _17623_/CLK _15828_/D vssd1 vssd1 vccd1 vccd1 _15828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15759_ _17680_/CLK _15759_/D vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08300_ hold1577/X _08336_/A2 _08299_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09280_ _12654_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _16251_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08231_ hold1190/X _08263_/A2 _08230_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08231_/X
+ sky130_fd_sc_hd__o211a_1
X_17429_ _17429_/CLK _17429_/D vssd1 vssd1 vccd1 vccd1 _17429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _15513_/A hold2506/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08093_ hold1241/X _08088_/B _08092_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4203 hold5893/X vssd1 vssd1 vccd1 vccd1 hold5894/A sky130_fd_sc_hd__buf_6
XFILLER_0_144_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4214 _13615_/X vssd1 vssd1 vccd1 vccd1 _17658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4225 _17687_/Q vssd1 vssd1 vccd1 vccd1 hold4225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4236 _12046_/X vssd1 vssd1 vccd1 vccd1 _17172_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4247 _17657_/Q vssd1 vssd1 vccd1 vccd1 hold4247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3502 _17279_/Q vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3513 hold5865/X vssd1 vssd1 vccd1 vccd1 hold5866/A sky130_fd_sc_hd__buf_6
Xhold4258 _12076_/X vssd1 vssd1 vccd1 vccd1 _17182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3524 _11407_/X vssd1 vssd1 vccd1 vccd1 _16959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4269 _17607_/Q vssd1 vssd1 vccd1 vccd1 hold4269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3535 _16844_/Q vssd1 vssd1 vccd1 vccd1 hold3535/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3546 _10599_/Y vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2801 _08024_/X vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2812 _18162_/Q vssd1 vssd1 vccd1 vccd1 hold2812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3557 _17358_/Q vssd1 vssd1 vccd1 vccd1 hold3557/X sky130_fd_sc_hd__dlygate4sd3_1
X_08995_ hold498/X _16115_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__mux2_1
XFILLER_0_228_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2823 _17982_/Q vssd1 vssd1 vccd1 vccd1 hold2823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3568 _11745_/Y vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2834 _17820_/Q vssd1 vssd1 vccd1 vccd1 hold2834/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3579 _16905_/Q vssd1 vssd1 vccd1 vccd1 hold3579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2845 _15538_/X vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07946_ _14116_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07946_/X sky130_fd_sc_hd__or2_1
Xhold2856 _17782_/Q vssd1 vssd1 vccd1 vccd1 hold2856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2867 _15838_/Q vssd1 vssd1 vccd1 vccd1 hold2867/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2878 _18156_/Q vssd1 vssd1 vccd1 vccd1 hold2878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2889 _13953_/X vssd1 vssd1 vccd1 vccd1 _17781_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07877_ _15555_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09616_ hold5387/X _11159_/B _09615_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _09616_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ hold3880/X _10007_/B _09546_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09547_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09478_ _09483_/C _09484_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _16320_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08429_ _14878_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ hold4038/X _11726_/B _11439_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ hold5581/X _11753_/B _11370_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11371_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ hold2339/X hold3744/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__mux2_1
X_13110_ _13110_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__or2_1
X_14090_ _15543_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _17522_/Q hold931/X _17523_/Q vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__or3b_1
Xhold5460 _13411_/X vssd1 vssd1 vccd1 vccd1 _17590_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10253_ hold1731/X _16575_/Q _10613_/C vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__mux2_1
Xhold5471 _16811_/Q vssd1 vssd1 vccd1 vccd1 hold5471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5482 _10753_/X vssd1 vssd1 vccd1 vccd1 _16741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5493 _16709_/Q vssd1 vssd1 vccd1 vccd1 hold5493/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4770 _09595_/X vssd1 vssd1 vccd1 vccd1 _16355_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10184_ hold2941/X _16552_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__mux2_1
Xhold4781 _16824_/Q vssd1 vssd1 vccd1 vccd1 hold4781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4792 _10102_/X vssd1 vssd1 vccd1 vccd1 _16524_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16800_ _18064_/CLK _16800_/D vssd1 vssd1 vccd1 vccd1 _16800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17780_ _17907_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_135_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14992_ _15099_/A _15016_/B vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout270 fanout334/X vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout281 _12273_/A vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__buf_4
X_16731_ _18050_/CLK _16731_/D vssd1 vssd1 vccd1 vccd1 _16731_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout292 _11124_/A vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13943_ _13943_/A _13943_/B vssd1 vssd1 vccd1 vccd1 _17777_/D sky130_fd_sc_hd__and2_1
XFILLER_0_221_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16662_ _18198_/CLK _16662_/D vssd1 vssd1 vccd1 vccd1 _16662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13874_ _17745_/Q _13886_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13874_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18401_ _18401_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15613_ _17145_/CLK _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _12912_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _17451_/D sky130_fd_sc_hd__and2_1
XFILLER_0_232_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16593_ _18181_/CLK _16593_/D vssd1 vssd1 vccd1 vccd1 _16593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _18364_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ hold2040/X _15560_/A2 _15543_/Y _15548_/C1 vssd1 vssd1 vccd1 vccd1 _15544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12756_ _12759_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _17428_/D sky130_fd_sc_hd__and2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18263_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ hold4463/X _11801_/B _11706_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11707_/X
+ sky130_fd_sc_hd__o211a_1
X_15475_ hold881/X _09386_/A _09362_/D hold776/X vssd1 vssd1 vccd1 vccd1 _15475_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ _12768_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _17405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17214_ _17234_/CLK _17214_/D vssd1 vssd1 vccd1 vccd1 _17214_/Q sky130_fd_sc_hd__dfxtp_1
X_14426_ hold3010/X _14433_/B _14425_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _14426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18194_ _18226_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ _11732_/A _11729_/B _11637_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _11638_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17145_ _17145_/CLK _17145_/D vssd1 vssd1 vccd1 vccd1 _17145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14357_ _14984_/A hold3099/X hold333/X vssd1 vssd1 vccd1 vccd1 _14358_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ hold5650/X _11789_/B _11568_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _11569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold707 hold707/A vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ hold4992/X _13307_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13308_/X sky130_fd_sc_hd__mux2_2
Xhold718 input53/X vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_208_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold729 la_data_in[29] vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ _17860_/CLK _17076_/D vssd1 vssd1 vccd1 vccd1 _17076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ _14968_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14288_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16027_ _16131_/CLK _16027_/D vssd1 vssd1 vccd1 vccd1 hold701/A sky130_fd_sc_hd__dfxtp_1
X_13239_ _13311_/A1 _13237_/X _13238_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2108 _08085_/X vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 _16234_/Q vssd1 vssd1 vccd1 vccd1 hold2119/X sky130_fd_sc_hd__dlygate4sd3_1
X_07800_ _18459_/Q _18457_/Q vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__nor2_1
X_08780_ _15414_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _16010_/D sky130_fd_sc_hd__and2_1
Xhold1407 _14444_/X vssd1 vssd1 vccd1 vccd1 _18018_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17978_ _18010_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1418 _15749_/Q vssd1 vssd1 vccd1 vccd1 hold1418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1429 _17765_/Q vssd1 vssd1 vccd1 vccd1 hold1429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16929_ _17871_/CLK _16929_/D vssd1 vssd1 vccd1 vccd1 _16929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _15231_/A _16286_/Q _09401_/S vssd1 vssd1 vccd1 vccd1 _09401_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_220_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09332_ hold1296/X _09338_/A2 _09331_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09263_ _15539_/A hold2531/X _09273_/S vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ hold2555/X _08213_/B _08213_/Y _08153_/A vssd1 vssd1 vccd1 vccd1 _08214_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ _15523_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08145_ _08145_/A _08145_/B vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _14529_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4000 _16401_/Q vssd1 vssd1 vccd1 vccd1 hold4000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4011 _13423_/X vssd1 vssd1 vccd1 vccd1 _17594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4022 _16630_/Q vssd1 vssd1 vccd1 vccd1 hold4022/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4033 _13426_/X vssd1 vssd1 vccd1 vccd1 _17595_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4044 _17628_/Q vssd1 vssd1 vccd1 vccd1 hold4044/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4055 _16887_/Q vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3310 _17384_/Q vssd1 vssd1 vccd1 vccd1 hold3310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4066 _10360_/X vssd1 vssd1 vccd1 vccd1 _16610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3321 _12369_/Y vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4077 _16465_/Q vssd1 vssd1 vccd1 vccd1 hold4077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3332 _12638_/X vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3343 _16652_/Q vssd1 vssd1 vccd1 vccd1 hold3343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4088 _11854_/X vssd1 vssd1 vccd1 vccd1 _17108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4099 _16679_/Q vssd1 vssd1 vccd1 vccd1 hold4099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3354 _12830_/X vssd1 vssd1 vccd1 vccd1 _12831_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3365 _16406_/Q vssd1 vssd1 vccd1 vccd1 hold3365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2620 _18039_/Q vssd1 vssd1 vccd1 vccd1 hold2620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkbuf_2
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3376 _09901_/X vssd1 vssd1 vccd1 vccd1 _16457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 _09105_/X vssd1 vssd1 vccd1 vccd1 _16167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3387 _09739_/X vssd1 vssd1 vccd1 vccd1 _16403_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2642 _17755_/Q vssd1 vssd1 vccd1 vccd1 hold2642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _13037_/A hold463/X vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__and2_1
XFILLER_0_215_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2653 _14637_/X vssd1 vssd1 vccd1 vccd1 _18109_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3398 _12842_/X vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__buf_4
Xhold2664 _17990_/Q vssd1 vssd1 vccd1 vccd1 hold2664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1930 _08432_/X vssd1 vssd1 vccd1 vccd1 _15846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 _08261_/X vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 _18149_/Q vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2686 _14959_/X vssd1 vssd1 vccd1 vccd1 _18264_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07929_ hold1159/X _07924_/B _07928_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _07929_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1952 _18157_/Q vssd1 vssd1 vccd1 vccd1 hold1952/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2697 _17808_/Q vssd1 vssd1 vccd1 vccd1 hold2697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 _14741_/X vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1974 _14181_/X vssd1 vssd1 vccd1 vccd1 _17891_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1985 _18328_/Q vssd1 vssd1 vccd1 vccd1 hold1985/X sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ hold1267/X _16804_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__mux2_1
Xhold1996 _18354_/Q vssd1 vssd1 vccd1 vccd1 hold1996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10871_ hold2823/X hold5178/X _11159_/C vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ hold1897/X hold3292/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13590_ _13791_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ hold1583/X _17358_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ hold324/X _15486_/A2 _09357_/B hold473/X vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a22o_1
X_12472_ _17329_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ hold2594/X _14198_/B _14210_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14211_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11423_ hold2306/X _16965_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__mux2_1
X_15191_ _15191_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14142_ _14946_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__nand2_1
X_11354_ hold3057/X hold5200/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11355_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_387_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17278_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ _10497_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14073_ hold1975/X _14107_/A2 _14072_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14073_/X
+ sky130_fd_sc_hd__o211a_1
X_11285_ hold1429/X hold5068/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_316_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18035_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5290 _17129_/Q vssd1 vssd1 vccd1 vccd1 hold5290/X sky130_fd_sc_hd__dlygate4sd3_1
X_13024_ hold990/X hold957/X vssd1 vssd1 vccd1 vccd1 _13025_/C sky130_fd_sc_hd__nand2_1
X_10236_ _10524_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__or2_1
X_17901_ _17901_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17832_ _17896_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10167_ _10527_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _18003_/CLK _17763_/D vssd1 vssd1 vccd1 vccd1 _17763_/Q sky130_fd_sc_hd__dfxtp_1
X_10098_ _10482_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14975_ hold1479/X hold514/X _14974_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16714_ _18429_/CLK _16714_/D vssd1 vssd1 vccd1 vccd1 _16714_/Q sky130_fd_sc_hd__dfxtp_1
X_13926_ hold469/X hold697/X hold124/X vssd1 vssd1 vccd1 vccd1 hold698/A sky130_fd_sc_hd__mux2_1
XFILLER_0_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17694_ _17694_/CLK _17694_/D vssd1 vssd1 vccd1 vccd1 _17694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16645_ _18201_/CLK _16645_/D vssd1 vssd1 vccd1 vccd1 _16645_/Q sky130_fd_sc_hd__dfxtp_1
X_13857_ hold3647/X _13776_/A _13856_/X vssd1 vssd1 vccd1 vccd1 _13857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12808_ hold1216/X hold3183/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16576_ _18164_/CLK _16576_/D vssd1 vssd1 vccd1 vccd1 _16576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13788_ _13788_/A _13788_/B vssd1 vssd1 vccd1 vccd1 _13788_/X sky130_fd_sc_hd__or2_1
X_18315_ _18321_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15527_ hold944/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15527_/X sky130_fd_sc_hd__or2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12739_ _16244_/Q _17424_/Q _12748_/S vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17879_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ _18366_/CLK hold928/X vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15458_ hold184/X _09367_/A _15479_/B1 _16022_/Q vssd1 vssd1 vccd1 vccd1 _15458_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14409_ _14517_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__or2_1
X_18177_ _18209_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
X_15389_ hold816/X _09365_/B _09392_/C hold901/X _15388_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _17160_/CLK _17128_/D vssd1 vssd1 vccd1 vccd1 _17128_/Q sky130_fd_sc_hd__dfxtp_1
Xhold515 hold515/A vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold526 hold526/A vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold537 hold537/A vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold548 hold548/A vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ hold1893/X hold4801/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__mux2_1
Xhold559 hold559/A vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__clkbuf_16
X_17059_ _17905_/CLK _17059_/D vssd1 vssd1 vccd1 vccd1 _17059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08901_ _15344_/A hold853/X vssd1 vssd1 vccd1 vccd1 _16068_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09881_ hold1204/X _16451_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ hold118/X hold610/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _18362_/Q vssd1 vssd1 vccd1 vccd1 hold1204/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _14891_/X vssd1 vssd1 vccd1 vccd1 _18232_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _08406_/X vssd1 vssd1 vccd1 vccd1 _15833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _18438_/Q vssd1 vssd1 vccd1 vccd1 hold1237/X sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ hold256/X _16002_/Q _08779_/S vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__mux2_1
Xhold1248 hold1277/X vssd1 vssd1 vccd1 vccd1 hold1248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1259 _08038_/X vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _15364_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _15968_/D sky130_fd_sc_hd__and2_1
XFILLER_0_196_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ _15103_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09246_ _12759_/A _09246_/B vssd1 vssd1 vccd1 vccd1 _16234_/D sky130_fd_sc_hd__and2_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09177_ hold1714/X _09177_/A2 _09176_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08128_ _15533_/A hold2864/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ hold2072/X _08097_/A2 _08058_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _08059_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11070_ _11070_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__or2_1
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput79 _13185_/A vssd1 vssd1 vccd1 vccd1 output79/X sky130_fd_sc_hd__buf_6
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3140 _15136_/X vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10021_ _11203_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _16497_/D sky130_fd_sc_hd__nor2_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3151 _18323_/Q vssd1 vssd1 vccd1 vccd1 hold3151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3162 _12905_/X vssd1 vssd1 vccd1 vccd1 _12906_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3173 _17473_/Q vssd1 vssd1 vccd1 vccd1 hold3173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3184 _17451_/Q vssd1 vssd1 vccd1 vccd1 hold3184/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3195 _17425_/Q vssd1 vssd1 vccd1 vccd1 hold3195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2450 _14335_/X vssd1 vssd1 vccd1 vccd1 _17965_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2461 _15865_/Q vssd1 vssd1 vccd1 vccd1 hold2461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 _08079_/X vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _08440_/X vssd1 vssd1 vccd1 vccd1 _15850_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2494 _17798_/Q vssd1 vssd1 vccd1 vccd1 hold2494/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1760 _14111_/X vssd1 vssd1 vccd1 vccd1 _17857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14760_ _15099_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__or2_1
Xhold1771 _18112_/Q vssd1 vssd1 vccd1 vccd1 hold1771/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1782 _14504_/X vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11972_ hold2384/X hold5443/X _13862_/C vssd1 vssd1 vccd1 vccd1 _11973_/B sky130_fd_sc_hd__mux2_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _15775_/Q vssd1 vssd1 vccd1 vccd1 hold1793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ hold3854/X _13814_/B _13710_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13711_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10923_ _11115_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__or2_1
X_14691_ hold2380/X _14720_/B _14690_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14691_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16430_ _18341_/CLK _16430_/D vssd1 vssd1 vccd1 vccd1 _16430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13642_ hold5727/X _13832_/B _13641_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13642_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _11052_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _18272_/CLK _16361_/D vssd1 vssd1 vccd1 vccd1 _16361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ hold4575/X _13847_/B _13572_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13573_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ _11070_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10785_/X sky130_fd_sc_hd__or2_1
X_18100_ _18164_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15312_ _15489_/A _15312_/B _15312_/C _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/X
+ sky130_fd_sc_hd__or4_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ hold3259/X _12523_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12524_/X sky130_fd_sc_hd__mux2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16312_/CLK _16292_/D vssd1 vssd1 vccd1 vccd1 _16292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _18063_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _15490_/A1 _15235_/X _15242_/X _15490_/B1 hold4271/X vssd1 vssd1 vccd1 vccd1
+ _15243_/X sky130_fd_sc_hd__a32o_1
X_12455_ hold88/X _12509_/A2 _12507_/A3 _12454_/X _12424_/A vssd1 vssd1 vccd1 vccd1
+ hold69/A sky130_fd_sc_hd__o311a_1
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ _12057_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15174_ hold5987/X _15165_/B hold1143/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _15174_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _12386_/A hold408/X vssd1 vssd1 vccd1 vccd1 _17286_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ hold1668/X _14142_/B _14124_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _14125_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11337_ _12204_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_150_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _14164_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11268_ _12219_/A _11268_/B vssd1 vssd1 vccd1 vccd1 _11268_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ hold999/X _13017_/B vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__or2_1
X_10219_ hold3944/X _10637_/B _10218_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11199_ hold4676/X _11103_/A _11198_/X vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17815_ _17815_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17746_ _17746_/CLK _17746_/D vssd1 vssd1 vccd1 vccd1 _17746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14958_ _15227_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13909_ _13909_/A _13909_/B vssd1 vssd1 vccd1 vccd1 _17760_/D sky130_fd_sc_hd__and2_1
X_17677_ _17677_/CLK _17677_/D vssd1 vssd1 vccd1 vccd1 _17677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14889_ hold2931/X _14880_/B _14888_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_43_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_43_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16628_ _18152_/CLK _16628_/D vssd1 vssd1 vccd1 vccd1 _16628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16559_ _18159_/CLK _16559_/D vssd1 vssd1 vccd1 vccd1 _16559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09100_ _15541_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ _12438_/A hold347/X vssd1 vssd1 vccd1 vccd1 _16132_/D sky130_fd_sc_hd__and2_1
X_18229_ _18229_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_238_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 hold334/A vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold345 input11/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__clkbuf_8
Xhold378 input13/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__or2_1
Xhold389 hold389/A vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout803 _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__buf_4
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 _15062_/A vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__buf_4
XFILLER_0_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout825 _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout836 _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ _09960_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__or2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 _07787_/Y vssd1 vssd1 vccd1 vccd1 fanout847/X sky130_fd_sc_hd__buf_8
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 _15221_/A vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__buf_12
Xhold1001 _18229_/Q vssd1 vssd1 vccd1 vccd1 hold1001/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 fanout873/X vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__buf_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1012 hold6043/X vssd1 vssd1 vccd1 vccd1 hold381/A sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _15491_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _16026_/D sky130_fd_sc_hd__and2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _15692_/Q vssd1 vssd1 vccd1 vccd1 hold1023/X sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _09963_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__or2_1
Xhold1034 hold1034/A vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 la_data_in[11] vssd1 vssd1 vccd1 vccd1 hold1045/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _17979_/Q vssd1 vssd1 vccd1 vccd1 hold1056/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 hold1067/A vssd1 vssd1 vccd1 vccd1 _15173_/A sky130_fd_sc_hd__clkbuf_16
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _15264_/A hold612/X vssd1 vssd1 vccd1 vccd1 _15993_/D sky130_fd_sc_hd__and2_1
Xhold1078 hold1154/X vssd1 vssd1 vccd1 vccd1 hold1155/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1089 _08508_/X vssd1 vssd1 vccd1 vccd1 _15881_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ hold47/X hold456/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__mux2_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _11194_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _16680_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ hold1680/X _09216_/B _09228_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _09229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _13461_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _12267_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11122_ hold5154/X _11216_/B _11121_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11122_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold890 hold890/A vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15930_ _17313_/CLK _15930_/D vssd1 vssd1 vccd1 vccd1 hold546/A sky130_fd_sc_hd__dfxtp_1
X_11053_ hold4489/X _11147_/B _11052_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _11053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _16492_/Q _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_1414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _17680_/CLK _15861_/D vssd1 vssd1 vccd1 vccd1 _15861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 _18087_/Q vssd1 vssd1 vccd1 vccd1 hold2280/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17696_/CLK _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2291 _18083_/Q vssd1 vssd1 vccd1 vccd1 hold2291/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _15205_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__or2_1
XFILLER_0_216_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _17723_/CLK _15792_/D vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _17534_/CLK _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1590 _14071_/X vssd1 vssd1 vccd1 vccd1 _17838_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14743_ hold3130/X _14774_/B _14742_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14743_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11955_ _12051_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ hold4781/X _11180_/B _10905_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10906_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17462_ _17482_/CLK _17462_/D vssd1 vssd1 vccd1 vccd1 _17462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14674_ _14782_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _12057_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16413_ _18292_/CLK _16413_/D vssd1 vssd1 vccd1 vccd1 _16413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ hold2085/X hold5685/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__mux2_1
X_17393_ _18442_/CLK _17393_/D vssd1 vssd1 vccd1 vccd1 _17393_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ hold4523/X _11789_/B _10836_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _10837_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ _18142_/CLK _16344_/D vssd1 vssd1 vccd1 vccd1 _16344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13556_ hold2264/X _17639_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ hold3894/X _11726_/B _10767_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _10768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12507_ hold77/X _08597_/Y _12507_/A3 _12506_/X _09053_/A vssd1 vssd1 vccd1 vccd1
+ hold78/A sky130_fd_sc_hd__o311a_1
XFILLER_0_171_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ _17517_/CLK _16275_/D vssd1 vssd1 vccd1 vccd1 _16275_/Q sky130_fd_sc_hd__dfxtp_1
X_13487_ hold1487/X _17616_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13488_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_331_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17872_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10699_ hold5016/X _11177_/B _10698_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__o211a_1
X_18014_ _18014_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ hold1470/X _15221_/B _15225_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _12438_/A hold168/X vssd1 vssd1 vccd1 vccd1 _17312_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15211_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15157_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12369_ hold3320/X _12273_/A _12368_/X vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3909 _10294_/X vssd1 vssd1 vccd1 vccd1 _16588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14108_ _14789_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_121_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15088_ hold1074/X _15111_/B _15087_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15088_/X
+ sky130_fd_sc_hd__o211a_1
X_14039_ hold1925/X _14038_/B _14038_/Y _13903_/A vssd1 vssd1 vccd1 vccd1 _14039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08600_ _12386_/A hold677/X vssd1 vssd1 vccd1 vccd1 _15922_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09580_ hold5669/X _10070_/B _09579_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09580_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08531_ _13046_/C _12380_/A vssd1 vssd1 vccd1 vccd1 _08536_/S sky130_fd_sc_hd__or2_2
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17729_ _17729_/CLK _17729_/D vssd1 vssd1 vccd1 vccd1 _17729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08462_ _14246_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08393_ hold203/X hold754/X vssd1 vssd1 vccd1 vccd1 _08393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_419_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17157_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ hold596/X _16124_/Q _09062_/S vssd1 vssd1 vccd1 vccd1 hold597/A sky130_fd_sc_hd__mux2_1
XFILLER_0_116_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5801 hold5938/X vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5812 output98/X vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_147_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5823 output97/X vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_12
Xhold5834 hold5834/A vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5845 _18406_/Q vssd1 vssd1 vccd1 vccd1 hold5845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold388/X vssd1 vssd1 vccd1 vccd1 hold389/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold763/X vssd1 vssd1 vccd1 vccd1 hold764/A sky130_fd_sc_hd__buf_4
Xhold5856 hold5856/A vssd1 vssd1 vccd1 vccd1 hold5856/X sky130_fd_sc_hd__clkbuf_4
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5867 hold6012/X vssd1 vssd1 vccd1 vccd1 hold5867/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold153 hold16/X vssd1 vssd1 vccd1 vccd1 input32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5878 hold5878/A vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_12
Xhold5889 _18411_/Q vssd1 vssd1 vccd1 vccd1 hold5889/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _12967_/S vssd1 vssd1 vccd1 vccd1 _12601_/S sky130_fd_sc_hd__buf_6
Xfanout611 _09362_/C vssd1 vssd1 vccd1 vccd1 _15479_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09916_ hold3886/X _10010_/B _09915_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09916_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout622 _15484_/A2 vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__buf_6
Xfanout633 _13304_/B1 vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__buf_6
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 fanout693/X vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__buf_2
Xfanout655 fanout693/X vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout666 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__buf_4
X_09847_ hold4739/X _10055_/B _09846_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout677 _08155_/A vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__buf_4
XFILLER_0_232_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 fanout692/X vssd1 vssd1 vccd1 vccd1 _14013_/C1 sky130_fd_sc_hd__buf_2
Xfanout699 _12386_/A vssd1 vssd1 vccd1 vccd1 _15264_/A sky130_fd_sc_hd__buf_4
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ hold4765/X _10049_/B _09777_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09778_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _17519_/Q _17518_/Q vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__nand2b_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11740_ _12310_/A _11740_/B vssd1 vssd1 vccd1 vccd1 _17070_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ hold5609/X _11789_/B _11670_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11671_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13410_ _13794_/A _13410_/B vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10622_ _16698_/Q _10622_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10622_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14390_ _14390_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _17992_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ _13698_/A _13341_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10553_ hold2931/X hold3776/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__mux2_1
X_16060_ _16322_/CLK _16060_/D vssd1 vssd1 vccd1 vccd1 hold889/A sky130_fd_sc_hd__dfxtp_1
X_13272_ _13265_/X _13271_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_121_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10484_ hold2778/X hold3343/X _10580_/C vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ hold1342/X _15004_/B _15010_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12223_ hold5258/X _12317_/B _12222_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _12223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12154_ hold3994/X _12374_/B _12153_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12154_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11105_ hold3104/X _16859_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12085_ hold4517/X _13877_/B _12084_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12085_/X
+ sky130_fd_sc_hd__o211a_1
X_16962_ _17904_/CLK _16962_/D vssd1 vssd1 vccd1 vccd1 _16962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15913_ _18407_/CLK _15913_/D vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__dfxtp_1
X_11036_ hold2075/X hold4119/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16893_ _17966_/CLK _16893_/D vssd1 vssd1 vccd1 vccd1 _16893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15844_ _17607_/CLK _15844_/D vssd1 vssd1 vccd1 vccd1 _15844_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _17694_/CLK _15775_/D vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12987_/A _12987_/B vssd1 vssd1 vccd1 vccd1 _17505_/D sky130_fd_sc_hd__and2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14726_ _14726_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__or2_1
X_17514_ _17515_/CLK _17514_/D vssd1 vssd1 vccd1 vccd1 _17514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11938_ hold5366/X _12353_/B _11937_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _11938_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17445_ _17446_/CLK _17445_/D vssd1 vssd1 vccd1 vccd1 _17445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ hold3051/X _14664_/B _14656_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11869_ hold4125/X _13868_/B _11868_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ _13800_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _17376_/CLK _17376_/D vssd1 vssd1 vccd1 vccd1 _17376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _15197_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14588_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16327_ _18272_/CLK _16327_/D vssd1 vssd1 vccd1 vccd1 _16327_/Q sky130_fd_sc_hd__dfxtp_1
X_13539_ _13767_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16258_ _17379_/CLK _16258_/D vssd1 vssd1 vccd1 vccd1 _16258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5108 _16783_/Q vssd1 vssd1 vccd1 vccd1 hold5108/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5119 _09892_/X vssd1 vssd1 vccd1 vccd1 _16454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _15209_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4407 _16743_/Q vssd1 vssd1 vccd1 vccd1 hold4407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16189_ _17877_/CLK _16189_/D vssd1 vssd1 vccd1 vccd1 _16189_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4418 _12151_/X vssd1 vssd1 vccd1 vccd1 _17207_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4429 _16894_/Q vssd1 vssd1 vccd1 vccd1 _11210_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3706 _17688_/Q vssd1 vssd1 vccd1 vccd1 hold3706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3717 _10291_/X vssd1 vssd1 vccd1 vccd1 _16587_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3728 _16575_/Q vssd1 vssd1 vccd1 vccd1 hold3728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3739 _13881_/Y vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07962_ _15531_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ hold3092/X _16391_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07893_ hold2586/X _07918_/B _07892_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09632_ hold1497/X _16368_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ hold1827/X _13230_/A _10481_/S vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_195_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ hold2056/X _08503_/Y _08513_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _08514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__or3_4
XFILLER_0_188_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08445_ _14894_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_253_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18228_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08376_ hold181/X _15820_/Q hold134/X vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5620 _11131_/X vssd1 vssd1 vccd1 vccd1 _16867_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5631 _16795_/Q vssd1 vssd1 vccd1 vccd1 hold5631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5642 _11665_/X vssd1 vssd1 vccd1 vccd1 _17045_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5653 _10041_/Y vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5664 _13827_/Y vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4930 _16597_/Q vssd1 vssd1 vccd1 vccd1 hold4930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5675 _16412_/Q vssd1 vssd1 vccd1 vccd1 hold5675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5686 _13531_/X vssd1 vssd1 vccd1 vccd1 _17630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4941 _12112_/X vssd1 vssd1 vccd1 vccd1 _17194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4952 _17110_/Q vssd1 vssd1 vccd1 vccd1 hold4952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5697 _17631_/Q vssd1 vssd1 vccd1 vccd1 hold5697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4963 _11208_/Y vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4974 _16639_/Q vssd1 vssd1 vccd1 vccd1 hold4974/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4985 _11754_/Y vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4996 _16965_/Q vssd1 vssd1 vccd1 vccd1 hold4996/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout430 _13311_/A1 vssd1 vssd1 vccd1 vccd1 _13199_/A1 sky130_fd_sc_hd__buf_8
Xfanout441 _12029_/S vssd1 vssd1 vccd1 vccd1 _13793_/S sky130_fd_sc_hd__clkbuf_8
Xfanout452 _11150_/C vssd1 vssd1 vccd1 vccd1 _11747_/C sky130_fd_sc_hd__clkbuf_4
Xfanout463 _10025_/C vssd1 vssd1 vccd1 vccd1 _12251_/S sky130_fd_sc_hd__buf_4
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout474 _11204_/C vssd1 vssd1 vccd1 vccd1 _11762_/C sky130_fd_sc_hd__clkbuf_8
Xfanout485 _09824_/S vssd1 vssd1 vccd1 vccd1 _11159_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout496 _11096_/S vssd1 vssd1 vccd1 vccd1 _11177_/C sky130_fd_sc_hd__clkbuf_8
X_12910_ hold1521/X hold3383/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _14556_/A hold1412/X _09120_/Y hold1750/X vssd1 vssd1 vccd1 vccd1 _13890_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ hold1680/X _17458_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ hold1947/X _15560_/A2 _15559_/X _12696_/A vssd1 vssd1 vccd1 vccd1 _15560_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12772_ hold1052/X hold3338/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__mux2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14511_ _15191_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14511_/X sky130_fd_sc_hd__or2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _17065_/Q _11726_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__and3_1
X_15491_ _15491_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__and2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17898_/CLK _17230_/D vssd1 vssd1 vccd1 vccd1 _17230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ hold2874/X _14446_/A2 _14441_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _14442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11654_ hold2907/X _17042_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10605_ hold4630/X _10554_/A _10604_/X vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17161_ _17161_/CLK _17161_/D vssd1 vssd1 vccd1 vccd1 _17161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ hold469/X hold645/X hold333/X vssd1 vssd1 vccd1 vccd1 hold646/A sky130_fd_sc_hd__mux2_1
XFILLER_0_182_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11585_ hold2795/X _17019_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _17335_/CLK _16112_/D vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__dfxtp_1
X_13324_ hold3424/X _13802_/B _13323_/X _13714_/C1 vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__o211a_1
X_10536_ _10536_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17092_ _17188_/CLK _17092_/D vssd1 vssd1 vccd1 vccd1 _17092_/Q sky130_fd_sc_hd__dfxtp_1
X_16043_ _16087_/CLK _16043_/D vssd1 vssd1 vccd1 vccd1 hold901/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _13311_/A1 _13253_/X _13254_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13255_/X
+ sky130_fd_sc_hd__o211a_1
X_10467_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ hold2590/X hold4940/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_237_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18046_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13186_ _17574_/Q _17108_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_237_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10554_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ hold1269/X hold4191/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__mux2_1
X_17994_ _17994_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
X_12068_ hold2645/X _17180_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _12069_/B sky130_fd_sc_hd__mux2_1
X_16945_ _17855_/CLK _16945_/D vssd1 vssd1 vccd1 vccd1 _16945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11019_ _11667_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16876_ _18045_/CLK _16876_/D vssd1 vssd1 vccd1 vccd1 _16876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _17642_/CLK _15827_/D vssd1 vssd1 vccd1 vccd1 _15827_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _17677_/CLK _15758_/D vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14709_ hold1765/X _14720_/B _14708_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14709_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15689_ _17170_/CLK _15689_/D vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08230_ _14164_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _17429_/CLK _17428_/D vssd1 vssd1 vccd1 vccd1 _17428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08161_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _15718_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _17379_/CLK _17359_/D vssd1 vssd1 vccd1 vccd1 _17359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08092_ _14330_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4204 _15413_/X vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4215 _16784_/Q vssd1 vssd1 vccd1 vccd1 hold4215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4226 _13606_/X vssd1 vssd1 vccd1 vccd1 _17655_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4237 _17432_/Q vssd1 vssd1 vccd1 vccd1 hold4237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4248 _13516_/X vssd1 vssd1 vccd1 vccd1 _17625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3503 _12271_/X vssd1 vssd1 vccd1 vccd1 _17247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3514 _09397_/X vssd1 vssd1 vccd1 vccd1 _16285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4259 _17713_/Q vssd1 vssd1 vccd1 vccd1 hold4259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3525 _16962_/Q vssd1 vssd1 vccd1 vccd1 hold3525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3536 _10966_/X vssd1 vssd1 vccd1 vccd1 _16812_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2802 _17830_/Q vssd1 vssd1 vccd1 vccd1 hold2802/X sky130_fd_sc_hd__dlygate4sd3_1
X_08994_ _12444_/A hold517/X vssd1 vssd1 vccd1 vccd1 _16114_/D sky130_fd_sc_hd__and2_1
Xhold3547 _16528_/Q vssd1 vssd1 vccd1 vccd1 hold3547/X sky130_fd_sc_hd__clkbuf_2
Xhold2813 _14747_/X vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3558 _12545_/X vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3569 _17098_/Q vssd1 vssd1 vccd1 vccd1 hold3569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 _15677_/Q vssd1 vssd1 vccd1 vccd1 hold2824/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2835 _14033_/X vssd1 vssd1 vccd1 vccd1 _17820_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07945_ hold2828/X _07991_/A2 _07944_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07945_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2846 _17999_/Q vssd1 vssd1 vccd1 vccd1 hold2846/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2857 _13955_/X vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_2_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold2868 _08416_/X vssd1 vssd1 vccd1 vccd1 _15838_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2879 _14733_/X vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07876_ hold2560/X _07869_/B _07875_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _11064_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_434_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17695_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09546_ _09936_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09477_/A _16319_/Q _09477_/C vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__and3_1
XFILLER_0_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08428_ hold2295/X _08433_/B _08427_/Y _08151_/A vssd1 vssd1 vccd1 vccd1 _08428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ _12750_/A hold950/X vssd1 vssd1 vccd1 vccd1 _15811_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11658_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ hold3793/X _10477_/A2 _10320_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5450 _11350_/X vssd1 vssd1 vccd1 vccd1 _16940_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13040_ input2/X input1/X hold930/X hold918/X vssd1 vssd1 vccd1 vccd1 _13040_/X sky130_fd_sc_hd__or4b_1
X_10252_ hold3920/X _11198_/B _10251_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5461 _17147_/Q vssd1 vssd1 vccd1 vccd1 hold5461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5472 _10867_/X vssd1 vssd1 vccd1 vccd1 _16779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5483 _16741_/Q vssd1 vssd1 vccd1 vccd1 hold5483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5494 _11137_/X vssd1 vssd1 vccd1 vccd1 _16869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4760 _09556_/X vssd1 vssd1 vccd1 vccd1 _16342_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10183_ hold4835/X _10571_/B _10182_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10183_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4771 _16852_/Q vssd1 vssd1 vccd1 vccd1 hold4771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4782 _10906_/X vssd1 vssd1 vccd1 vccd1 _16792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4793 _16916_/Q vssd1 vssd1 vccd1 vccd1 hold4793/X sky130_fd_sc_hd__dlygate4sd3_1
X_14991_ hold1497/X hold514/X _14990_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _14991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout260 _11712_/A vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__buf_4
Xfanout271 _13776_/A vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__buf_4
Xfanout282 fanout334/X vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16730_ _18055_/CLK _16730_/D vssd1 vssd1 vccd1 vccd1 _16730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13942_ _14443_/A hold1234/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__mux2_1
Xfanout293 _11124_/A vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__buf_4
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16661_ _18219_/CLK _16661_/D vssd1 vssd1 vccd1 vccd1 _16661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _17744_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_175_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18389_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18400_ _18415_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_15612_ _17260_/CLK _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ hold3184/X _12823_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__mux2_1
X_16592_ _18186_/CLK _16592_/D vssd1 vssd1 vccd1 vccd1 _16592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18331_ _18331_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
X_15543_ _15543_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ hold3403/X _12754_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__mux2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18262_/CLK hold985/X vssd1 vssd1 vccd1 vccd1 hold984/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A _11706_/B vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__or2_1
X_15474_ hold176/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12686_ hold4168/X _12685_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__mux2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _15105_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14425_/X sky130_fd_sc_hd__or2_1
X_17213_ _17245_/CLK _17213_/D vssd1 vssd1 vccd1 vccd1 _17213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18193_ _18193_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17144_ _17872_/CLK _17144_/D vssd1 vssd1 vccd1 vccd1 _17144_/Q sky130_fd_sc_hd__dfxtp_1
X_14356_ _14356_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _17975_/D sky130_fd_sc_hd__and2_1
XFILLER_0_208_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11568_ _11670_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold708 hold708/A vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13307_ _13306_/X _16931_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__mux2_1
X_10519_ hold4942/X _10637_/B _10518_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10519_/X
+ sky130_fd_sc_hd__o211a_1
Xhold719 hold719/A vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__buf_8
X_17075_ _17825_/CLK _17075_/D vssd1 vssd1 vccd1 vccd1 _17075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14287_ hold754/X _14502_/B vssd1 vssd1 vccd1 vccd1 _14338_/B sky130_fd_sc_hd__or2_4
XFILLER_0_208_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _12234_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _18423_/CLK _16026_/D vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _13238_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13169_ _13169_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__and2_1
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2109 _18077_/Q vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ _18041_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1408 _17786_/Q vssd1 vssd1 vccd1 vccd1 hold1408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _08226_/X vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16928_ _17870_/CLK _16928_/D vssd1 vssd1 vccd1 vccd1 _16928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859_ _18060_/CLK _16859_/D vssd1 vssd1 vccd1 vccd1 _16859_/Q sky130_fd_sc_hd__dfxtp_1
X_09400_ _09400_/A _09400_/B _09400_/C vssd1 vssd1 vccd1 vccd1 _09401_/S sky130_fd_sc_hd__or3_1
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _15173_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09331_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _12738_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _16242_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08213_ _14774_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ hold2138/X _09218_/B _09192_/X _12807_/A vssd1 vssd1 vccd1 vccd1 _09193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _15549_/A hold2220/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08145_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08075_ hold2824/X _08097_/A2 _08074_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _08075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4001 _09637_/X vssd1 vssd1 vccd1 vccd1 _16369_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4012 _17582_/Q vssd1 vssd1 vccd1 vccd1 hold4012/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4023 _10324_/X vssd1 vssd1 vccd1 vccd1 _16598_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4034 _16459_/Q vssd1 vssd1 vccd1 vccd1 hold4034/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3300 _17372_/Q vssd1 vssd1 vccd1 vccd1 hold3300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4045 _13429_/X vssd1 vssd1 vccd1 vccd1 _17596_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3311 _12623_/X vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4056 _11095_/X vssd1 vssd1 vccd1 vccd1 _16855_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4067 _16580_/Q vssd1 vssd1 vccd1 vccd1 hold4067/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3322 _17483_/Q vssd1 vssd1 vccd1 vccd1 hold3322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4078 _09829_/X vssd1 vssd1 vccd1 vccd1 _16433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3333 _17445_/Q vssd1 vssd1 vccd1 vccd1 hold3333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3344 _10390_/X vssd1 vssd1 vccd1 vccd1 _16620_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4089 _17719_/Q vssd1 vssd1 vccd1 vccd1 hold4089/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2610 _08332_/X vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3355 _17455_/Q vssd1 vssd1 vccd1 vccd1 hold3355/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3366 _09652_/X vssd1 vssd1 vccd1 vccd1 _16374_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 _14488_/X vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08977_ hold228/X hold462/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__mux2_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2632 _18453_/Q vssd1 vssd1 vccd1 vccd1 hold2632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3377 _17475_/Q vssd1 vssd1 vccd1 vccd1 hold3377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__buf_4
Xhold3388 _16423_/Q vssd1 vssd1 vccd1 vccd1 hold3388/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2643 _15857_/Q vssd1 vssd1 vccd1 vccd1 hold2643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3399 _16393_/Q vssd1 vssd1 vccd1 vccd1 hold3399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 _18290_/Q vssd1 vssd1 vccd1 vccd1 hold2654/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1920 _09119_/X vssd1 vssd1 vccd1 vccd1 _16174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2665 _16214_/Q vssd1 vssd1 vccd1 vccd1 hold2665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 _18309_/Q vssd1 vssd1 vccd1 vccd1 hold2676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 _18170_/Q vssd1 vssd1 vccd1 vccd1 hold1931/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07928_ _15551_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07928_/X sky130_fd_sc_hd__or2_1
Xhold68 hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__clkbuf_2
Xhold1942 _14719_/X vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 _18124_/Q vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _14737_/X vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _14009_/X vssd1 vssd1 vccd1 vccd1 _17808_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 _18138_/Q vssd1 vssd1 vccd1 vccd1 hold1964/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1975 _17839_/Q vssd1 vssd1 vccd1 vccd1 hold1975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1986 _15092_/X vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _15537_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07859_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1997 _15146_/X vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10870_ hold5491/X _11156_/B _10869_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10870_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ hold3426/X _10025_/B _09528_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09529_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12606_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _17356_/D sky130_fd_sc_hd__and2_1
XFILLER_0_17_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ hold29/X _12445_/A _12445_/B _12470_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold30/A sky130_fd_sc_hd__o311a_1
XFILLER_0_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _15555_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11422_ hold3930/X _11747_/B _11421_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _11422_/X
+ sky130_fd_sc_hd__o211a_1
X_15190_ hold3201/X _15221_/B _15189_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14141_ hold1557/X _14142_/B _14140_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14141_/X
+ sky130_fd_sc_hd__o211a_1
X_11353_ hold5377/X _11732_/B _11352_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10304_ hold2172/X hold3742/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14072_ _15199_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11284_ hold5495/X _11762_/B _11283_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ hold990/X hold957/A vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__or2_1
Xhold5280 _16484_/Q vssd1 vssd1 vccd1 vccd1 hold5280/X sky130_fd_sc_hd__dlygate4sd3_1
X_17900_ _17900_/CLK _17900_/D vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_1
X_10235_ hold2532/X _16569_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5291 _11821_/X vssd1 vssd1 vccd1 vccd1 _17097_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4590 _09377_/X vssd1 vssd1 vccd1 vccd1 _16280_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17831_ _17863_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10166_ hold2371/X hold3607/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_206_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_356_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_234_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17762_ _17860_/CLK _17762_/D vssd1 vssd1 vccd1 vccd1 _17762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10097_ hold1865/X _16523_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__mux2_1
X_14974_ _14974_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_234_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ _18012_/CLK _16713_/D vssd1 vssd1 vccd1 vccd1 _16713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13925_ _13941_/A _13925_/B vssd1 vssd1 vccd1 vccd1 _17768_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17693_ _17693_/CLK _17693_/D vssd1 vssd1 vccd1 vccd1 _17693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_6_33_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_33_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ _18232_/CLK _16644_/D vssd1 vssd1 vccd1 vccd1 _16644_/Q sky130_fd_sc_hd__dfxtp_1
X_13856_ _17739_/Q _13856_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12807_ _12807_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _17445_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16575_ _18131_/CLK _16575_/D vssd1 vssd1 vccd1 vccd1 _16575_/Q sky130_fd_sc_hd__dfxtp_1
X_13787_ hold1414/X hold4197/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13788_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10999_ hold3914/X _11095_/A2 _10998_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18314_ _18346_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12738_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _17422_/D sky130_fd_sc_hd__and2_1
X_15526_ hold3023/X _15547_/B _15525_/X _12759_/A vssd1 vssd1 vccd1 vccd1 _15526_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15457_ hold799/X _09392_/C _15484_/B1 hold840/X _15456_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/B sky130_fd_sc_hd__a221o_1
X_18245_ _18379_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _12810_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _17399_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14408_ hold2681/X _14446_/A2 _14407_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ hold909/X _09386_/A _09392_/D hold795/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__a22o_1
X_18176_ _18176_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17127_ _17221_/CLK _17127_/D vssd1 vssd1 vccd1 vccd1 _17127_/Q sky130_fd_sc_hd__dfxtp_1
X_14339_ hold2899/X _14326_/B _14338_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14339_/X
+ sky130_fd_sc_hd__o211a_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold516 hold516/A vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 hold527/A vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold538 hold538/A vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _17904_/CLK _17058_/D vssd1 vssd1 vccd1 vccd1 _17058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 hold549/A vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16009_ _18422_/CLK _16009_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
X_08900_ hold346/X hold852/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__mux2_1
X_09880_ hold5094/X _10070_/B _09879_/X _09976_/C1 vssd1 vssd1 vccd1 vccd1 _09880_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _15304_/A hold863/X vssd1 vssd1 vccd1 vccd1 _16034_/D sky130_fd_sc_hd__and2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _15162_/X vssd1 vssd1 vccd1 vccd1 _18362_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1216 _16215_/Q vssd1 vssd1 vccd1 vccd1 hold1216/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _15324_/A hold728/X vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__and2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _16177_/Q vssd1 vssd1 vccd1 vccd1 hold1227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1238 _15524_/X vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1249 hold1249/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__buf_12
XFILLER_0_206_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08693_ hold118/X hold430/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ hold1779/X _09325_/B _09313_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _15521_/A hold2119/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09176_ _15559_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08127_ _08127_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08058_ _15517_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3130 _18160_/Q vssd1 vssd1 vccd1 vccd1 hold3130/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10020_ _13166_/A _11061_/A _10019_/X vssd1 vssd1 vccd1 vccd1 _10020_/Y sky130_fd_sc_hd__a21oi_1
Xhold3141 _18139_/Q vssd1 vssd1 vccd1 vccd1 hold3141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3152 _15082_/X vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3163 _17751_/Q vssd1 vssd1 vccd1 vccd1 hold3163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3174 _12890_/X vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3185 _17919_/Q vssd1 vssd1 vccd1 vccd1 hold3185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2440 _08497_/X vssd1 vssd1 vccd1 vccd1 _15877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2451 _15794_/Q vssd1 vssd1 vccd1 vccd1 hold2451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3196 _12746_/X vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2462 _08473_/X vssd1 vssd1 vccd1 vccd1 _15865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2473 _15602_/Q vssd1 vssd1 vccd1 vccd1 hold2473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 _18090_/Q vssd1 vssd1 vccd1 vccd1 hold2484/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1750 _13889_/Y vssd1 vssd1 vccd1 vccd1 hold1750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2495 _13987_/X vssd1 vssd1 vccd1 vccd1 _17798_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 _15641_/Q vssd1 vssd1 vccd1 vccd1 hold1761/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ hold5431/X _12353_/B _11970_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11971_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1772 _14643_/X vssd1 vssd1 vccd1 vccd1 _18112_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _17807_/Q vssd1 vssd1 vccd1 vccd1 hold1783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 _08281_/X vssd1 vssd1 vccd1 vccd1 _15775_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13710_ _13800_/A _13710_/B vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ hold2846/X _16798_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__mux2_1
X_14690_ _15191_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__or2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13641_ _13698_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _13641_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ hold3099/X _16775_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _18303_/CLK _16360_/D vssd1 vssd1 vccd1 vccd1 _16360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13746_/A _13572_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__or2_1
X_10784_ hold1281/X _16752_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__mux2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _09418_/B _09362_/A _15487_/B1 hold897/X _15310_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_137_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _17514_/Q _17352_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__mux2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16312_/CLK _16291_/D vssd1 vssd1 vccd1 vccd1 _16291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15242_ _15489_/A _15242_/B _15242_/C _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_164_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18030_ _18030_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_12454_ _17320_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ hold1704/X _16959_/Q _11480_/S vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__mux2_1
X_15173_ _15173_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12385_ hold215/X hold407/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold408/A sky130_fd_sc_hd__mux2_1
XFILLER_0_240_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _14517_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14124_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11336_ hold2856/X hold3928/X _11711_/S vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _14735_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__or2_4
X_11267_ hold2169/X hold3583/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ hold1716/X _13003_/Y _13005_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _13006_/X
+ sky130_fd_sc_hd__o211a_1
X_10218_ _10542_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11198_ _16890_/Q _11198_/B _11198_/C vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__and3_1
XTAP_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_190_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17814_ _17814_/CLK hold994/X vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__dfxtp_1
XTAP_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10149_ _10497_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17745_ _17745_/CLK _17745_/D vssd1 vssd1 vccd1 vccd1 _17745_/Q sky130_fd_sc_hd__dfxtp_1
X_14957_ hold1430/X _14952_/B _14956_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _14517_/A hold1507/X hold124/X vssd1 vssd1 vccd1 vccd1 _13908_/X sky130_fd_sc_hd__mux2_1
X_17676_ _17740_/CLK _17676_/D vssd1 vssd1 vccd1 vccd1 _17676_/Q sky130_fd_sc_hd__dfxtp_1
X_14888_ _15227_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16627_ _18215_/CLK _16627_/D vssd1 vssd1 vccd1 vccd1 _16627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13839_ _17573_/Q _13761_/A _13838_/X vssd1 vssd1 vccd1 vccd1 _13839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16558_ _18178_/CLK _16558_/D vssd1 vssd1 vccd1 vccd1 _16558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _15509_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16489_ _18367_/CLK _16489_/D vssd1 vssd1 vccd1 vccd1 _16489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ hold346/X _16132_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold347/A sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18228_ _18228_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18159_ _18159_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold346 hold41/X vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__buf_4
XFILLER_0_229_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_278_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18142_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09932_ hold1481/X hold3876/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__mux2_1
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold379 hold53/X vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_207_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18294_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout804 _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14392_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout815 _15026_/A vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout826 _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14797_/C1 sky130_fd_sc_hd__buf_4
X_09863_ hold1571/X _16445_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__mux2_1
Xfanout837 fanout847/X vssd1 vssd1 vccd1 vccd1 _14827_/C1 sky130_fd_sc_hd__buf_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout848 _07785_/Y vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__clkbuf_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 _07780_/Y vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__clkbuf_16
X_08814_ hold17/X hold433/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__mux2_1
Xhold1002 _14885_/X vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 hold381/X vssd1 vssd1 vccd1 vccd1 input41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 hold5839/X vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__clkbuf_4
X_09794_ _18333_/Q _16422_/Q _10034_/C vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__mux2_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1035 input65/X vssd1 vssd1 vccd1 vccd1 hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 hold1046/A vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ hold596/X hold611/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold612/A sky130_fd_sc_hd__mux2_1
Xhold1057 _16181_/Q vssd1 vssd1 vccd1 vccd1 hold1057/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 _14439_/X vssd1 vssd1 vccd1 vccd1 hold1068/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 hold1156/X vssd1 vssd1 vccd1 vccd1 hold1079/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _09015_/A _08676_/B vssd1 vssd1 vccd1 vccd1 _15959_/D sky130_fd_sc_hd__and2_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ _15557_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09159_ hold2395/X _09164_/B _09158_/Y _12894_/A vssd1 vssd1 vccd1 vccd1 _09159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ hold2422/X hold4257/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold880 hold880/A vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold891 hold891/A vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__or2_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10003_ _11203_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _16491_/D sky130_fd_sc_hd__nor2_1
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _17276_/CLK _15860_/D vssd1 vssd1 vccd1 vccd1 _15860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 _07979_/X vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2281 _14591_/X vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14811_ hold3025/X _14826_/B _14810_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14811_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2292 _14583_/X vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _17658_/CLK _15791_/D vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1580 _14823_/X vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17534_/CLK _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14742_ _15189_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__or2_1
Xhold1591 _18243_/Q vssd1 vssd1 vccd1 vccd1 hold1591/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11954_ hold2107/X _17142_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10905_ _11100_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__or2_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14673_ hold2774/X _14666_/B _14672_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14673_/X
+ sky130_fd_sc_hd__o211a_1
X_17461_ _17482_/CLK _17461_/D vssd1 vssd1 vccd1 vccd1 _17461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ hold2220/X hold3734/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16412_ _18323_/CLK _16412_/D vssd1 vssd1 vccd1 vccd1 _16412_/Q sky130_fd_sc_hd__dfxtp_1
X_13624_ hold3395/X _13808_/B _13623_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ _11670_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ _18442_/CLK _17392_/D vssd1 vssd1 vccd1 vccd1 _17392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16343_ _18390_/CLK _16343_/D vssd1 vssd1 vccd1 vccd1 _16343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13555_ hold4395/X _13847_/B _13554_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ _11631_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _17346_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16274_ _17376_/CLK _16274_/D vssd1 vssd1 vccd1 vccd1 _16274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ hold3517/X _13777_/A2 _13485_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _13486_/X
+ sky130_fd_sc_hd__o211a_1
X_10698_ _11082_/A _10698_/B vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15225_ _15225_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__or2_1
X_18013_ _18044_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12437_ hold140/X hold167/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__mux2_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15156_ hold1885/X _15167_/B _15155_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15156_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12368_ _17280_/Q _13877_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_371_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17701_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14107_ hold3012/X _14107_/A2 _14106_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ _11679_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__or2_1
X_15087_ _15195_/A hold734/X vssd1 vssd1 vccd1 vccd1 _15087_/X sky130_fd_sc_hd__or2_1
X_12299_ _17257_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_300_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17863_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14038_ _15004_/A _14038_/B vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15989_ _17304_/CLK _15989_/D vssd1 vssd1 vccd1 vccd1 hold767/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08530_ _13056_/C _17520_/Q _08868_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__or3_1
XFILLER_0_145_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17728_ _17728_/CLK _17728_/D vssd1 vssd1 vccd1 vccd1 _17728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08461_ hold1138/X _08488_/B _08460_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17659_ _17723_/CLK _17659_/D vssd1 vssd1 vccd1 vccd1 _17659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08392_ hold752/A hold689/A hold732/X hold764/A vssd1 vssd1 vccd1 vccd1 hold753/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_459_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09013_ _09063_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _16123_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5802 output82/X vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5813 hold5946/X vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__buf_1
XFILLER_0_182_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5824 hold5948/X vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__buf_1
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5835 _18408_/Q vssd1 vssd1 vccd1 vccd1 hold5835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold390/X vssd1 vssd1 vccd1 vccd1 hold391/A sky130_fd_sc_hd__buf_4
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold132 hold330/X vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_83_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5846 hold5846/A vssd1 vssd1 vccd1 vccd1 hold5846/X sky130_fd_sc_hd__buf_2
Xhold5857 _16280_/Q vssd1 vssd1 vccd1 vccd1 hold5857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold4/X vssd1 vssd1 vccd1 vccd1 input24/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5868 hold5868/A vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_12
Xhold154 input32/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5879 hold6015/X vssd1 vssd1 vccd1 vccd1 hold5879/X sky130_fd_sc_hd__buf_2
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _12970_/S vssd1 vssd1 vccd1 vccd1 _12967_/S sky130_fd_sc_hd__clkbuf_4
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _09358_/Y vssd1 vssd1 vccd1 vccd1 _15487_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_10_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09915_ _09933_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout623 _09347_/Y vssd1 vssd1 vccd1 vccd1 _15484_/A2 sky130_fd_sc_hd__buf_8
Xfanout634 _13304_/B1 vssd1 vssd1 vccd1 vccd1 _13312_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout645 _13714_/C1 vssd1 vssd1 vccd1 vccd1 _12738_/A sky130_fd_sc_hd__clkbuf_4
Xfanout656 _12987_/A vssd1 vssd1 vccd1 vccd1 _12996_/A sky130_fd_sc_hd__buf_4
X_09846_ _09960_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__or2_1
Xfanout667 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13720_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout678 _08155_/A vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__buf_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _14442_/C1 vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__buf_4
XFILLER_0_241_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09954_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _09015_/A hold151/X vssd1 vssd1 vccd1 vccd1 _15985_/D sky130_fd_sc_hd__and2_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ hold498/X hold909/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold910/A sky130_fd_sc_hd__mux2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__or2_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ _18461_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _16697_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13340_ hold2672/X hold5659/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ hold4075/X _10646_/B _10551_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13271_ _13311_/A1 _13269_/X _13270_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13271_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_126_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ _10577_/A _10577_/B _10482_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_129_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17303_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15010_ _15225_/A _15016_/B vssd1 vssd1 vccd1 vccd1 _15010_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _12285_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__or2_1
X_12153_ _13461_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ hold5164/X _11198_/B _11103_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _11104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12084_ _13782_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__or2_1
X_16961_ _17871_/CLK _16961_/D vssd1 vssd1 vccd1 vccd1 _16961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15912_ _18401_/CLK _15912_/D vssd1 vssd1 vccd1 vccd1 hold695/A sky130_fd_sc_hd__dfxtp_1
X_11035_ hold5286/X _11216_/B _11034_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16892_ _18061_/CLK _16892_/D vssd1 vssd1 vccd1 vccd1 _16892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _17702_/CLK _15843_/D vssd1 vssd1 vccd1 vccd1 _15843_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _17693_/CLK _15774_/D vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfxtp_1
X_12986_ hold3136/X _12985_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__mux2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17513_ _18398_/CLK _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ hold1569/X _14714_/B _14724_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14725_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _13794_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/CLK _17444_/D vssd1 vssd1 vccd1 vccd1 _17444_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _15103_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11868_ _13773_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10819_ hold5631/X _11201_/B _10818_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o211a_1
X_13607_ hold1462/X _17656_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__mux2_1
X_17375_ _17517_/CLK _17375_/D vssd1 vssd1 vccd1 vccd1 _17375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14587_ hold2397/X _14610_/B _14586_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14587_/X
+ sky130_fd_sc_hd__o211a_1
X_11799_ hold3852/X _12057_/A _11798_/X vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16326_ _18237_/CLK _16326_/D vssd1 vssd1 vccd1 vccd1 _16326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13538_ _15818_/Q _17633_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ _17379_/CLK _16257_/D vssd1 vssd1 vccd1 vccd1 _16257_/Q sky130_fd_sc_hd__dfxtp_1
X_13469_ hold2588/X hold3504/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13470_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5109 _10783_/X vssd1 vssd1 vccd1 vccd1 _16751_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15208_ hold1452/X _15219_/B _15207_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15208_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4408 _10663_/X vssd1 vssd1 vccd1 vccd1 _16711_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16188_ _17879_/CLK _16188_/D vssd1 vssd1 vccd1 vccd1 _16188_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4419 _16794_/Q vssd1 vssd1 vccd1 vccd1 hold4419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15139_ _15193_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15139_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3707 _13609_/X vssd1 vssd1 vccd1 vccd1 _17656_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3718 _16604_/Q vssd1 vssd1 vccd1 vccd1 hold3718/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3729 _10159_/X vssd1 vssd1 vccd1 vccd1 _16543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07961_ hold2905/X _07991_/A2 _07960_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07961_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09700_ hold5048/X _10034_/B _09699_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09700_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07892_ _14116_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09631_ hold3392/X _10010_/B _09630_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09631_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ hold5671/X _11177_/B _09561_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _09562_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08513_ _15517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 _09493_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_136_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08444_ hold1206/X _08433_/B _08443_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _12747_/A hold135/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_293_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17997_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_222_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18175_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5610 _11671_/X vssd1 vssd1 vccd1 vccd1 _17047_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5621 _16402_/Q vssd1 vssd1 vccd1 vccd1 hold5621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5632 _10819_/X vssd1 vssd1 vccd1 vccd1 _16763_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5643 _16866_/Q vssd1 vssd1 vccd1 vccd1 hold5643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5654 _16348_/Q vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4920 _11223_/Y vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5665 _16586_/Q vssd1 vssd1 vccd1 vccd1 hold5665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4931 _10225_/X vssd1 vssd1 vccd1 vccd1 _16565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5676 _09670_/X vssd1 vssd1 vccd1 vccd1 _16380_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4942 _16695_/Q vssd1 vssd1 vccd1 vccd1 hold4942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5687 _16548_/Q vssd1 vssd1 vccd1 vccd1 hold5687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5698 _13438_/X vssd1 vssd1 vccd1 vccd1 _17599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4953 _12339_/Y vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4964 _17092_/Q vssd1 vssd1 vccd1 vccd1 hold4964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4975 _10351_/X vssd1 vssd1 vccd1 vccd1 _16607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4986 _16671_/Q vssd1 vssd1 vccd1 vccd1 hold4986/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout420 _14000_/Y vssd1 vssd1 vccd1 vccd1 _14038_/B sky130_fd_sc_hd__buf_6
Xfanout431 _13052_/X vssd1 vssd1 vccd1 vccd1 _13311_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_195_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4997 _11329_/X vssd1 vssd1 vccd1 vccd1 _16933_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout442 _12029_/S vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__clkbuf_8
Xfanout453 _11168_/C vssd1 vssd1 vccd1 vccd1 _11732_/C sky130_fd_sc_hd__buf_6
Xfanout464 _13874_/C vssd1 vssd1 vccd1 vccd1 _13883_/C sky130_fd_sc_hd__clkbuf_8
Xfanout475 _11480_/S vssd1 vssd1 vccd1 vccd1 _11204_/C sky130_fd_sc_hd__buf_4
XFILLER_0_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout486 _09824_/S vssd1 vssd1 vccd1 vccd1 _11201_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_214_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09829_ hold4077/X _10010_/B _09828_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09829_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout497 _10580_/C vssd1 vssd1 vccd1 vccd1 _10190_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12870_/A _12840_/B vssd1 vssd1 vccd1 vccd1 _17456_/D sky130_fd_sc_hd__and2_1
XFILLER_0_214_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12780_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _17433_/D sky130_fd_sc_hd__and2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ hold1644/X _14535_/B _14509_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _14510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _12310_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _17064_/D sky130_fd_sc_hd__nor2_1
X_15490_ _15490_/A1 _15483_/X _15489_/X _15490_/B1 hold5896/A vssd1 vssd1 vccd1 vccd1
+ _15490_/X sky130_fd_sc_hd__a32o_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ hold3940/X _11747_/B _11652_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11653_/X
+ sky130_fd_sc_hd__o211a_1
X_14441_ _15229_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14441_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _16692_/Q _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__and3_1
X_14372_ _15032_/A _14372_/B vssd1 vssd1 vccd1 vccd1 _17983_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17160_ _17160_/CLK _17160_/D vssd1 vssd1 vccd1 vccd1 _17160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11584_ hold5547/X _11584_/A2 _11583_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16111_ _17334_/CLK _16111_/D vssd1 vssd1 vccd1 vccd1 hold436/A sky130_fd_sc_hd__dfxtp_1
X_13323_ _13800_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ hold1174/X _16669_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17091_ _17777_/CLK _17091_/D vssd1 vssd1 vccd1 vccd1 _17091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _17298_/CLK _16042_/D vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__dfxtp_1
X_13254_ _13254_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ hold1607/X _16646_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ hold5132/X _12299_/B _12204_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _12205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13185_ _13185_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__and2_1
XFILLER_0_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ hold2915/X _16623_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12136_ hold4229/X _13871_/B _12135_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17993_ _18053_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12067_ hold5435/X _12353_/B _12066_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o211a_1
X_16944_ _17851_/CLK _16944_/D vssd1 vssd1 vccd1 vccd1 _16944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18401_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11018_ hold2634/X hold4380/X _11204_/C vssd1 vssd1 vccd1 vccd1 _11019_/B sky130_fd_sc_hd__mux2_1
X_16875_ _18044_/CLK _16875_/D vssd1 vssd1 vccd1 vccd1 _16875_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15826_ _17641_/CLK _15826_/D vssd1 vssd1 vccd1 vccd1 _15826_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15757_ _17612_/CLK _15757_/D vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12969_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _17499_/D sky130_fd_sc_hd__and2_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ _15209_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14708_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ _17234_/CLK _15688_/D vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17427_ _17429_/CLK _17427_/D vssd1 vssd1 vccd1 vccd1 _17427_/Q sky130_fd_sc_hd__dfxtp_1
X_14639_ hold3063/X _14666_/B _14638_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08160_ hold999/X _15718_/Q _08170_/S vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__mux2_1
X_17358_ _17378_/CLK _17358_/D vssd1 vssd1 vccd1 vccd1 _17358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ _16312_/CLK _16309_/D vssd1 vssd1 vccd1 vccd1 _16309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ hold2210/X _08088_/B _08090_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08091_/X
+ sky130_fd_sc_hd__o211a_1
X_17289_ _18403_/CLK _17289_/D vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4205 _17197_/Q vssd1 vssd1 vccd1 vccd1 hold4205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4216 _10786_/X vssd1 vssd1 vccd1 vccd1 _16752_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4227 _17035_/Q vssd1 vssd1 vccd1 vccd1 hold4227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4238 _16746_/Q vssd1 vssd1 vccd1 vccd1 hold4238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4249 hold5835/X vssd1 vssd1 vccd1 vccd1 hold5836/A sky130_fd_sc_hd__buf_4
Xhold3504 _17610_/Q vssd1 vssd1 vccd1 vccd1 hold3504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3515 _16779_/Q vssd1 vssd1 vccd1 vccd1 hold3515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3526 _11320_/X vssd1 vssd1 vccd1 vccd1 _16930_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08993_ hold292/X hold516/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__mux2_1
Xhold3537 _16345_/Q vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_228_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3548 _10593_/Y vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2803 _14053_/X vssd1 vssd1 vccd1 vccd1 _17830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3559 _16334_/Q vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 _18043_/Q vssd1 vssd1 vccd1 vccd1 hold2814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 _08075_/X vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07944_ _15513_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07944_/X sky130_fd_sc_hd__or2_1
Xhold2836 _15788_/Q vssd1 vssd1 vccd1 vccd1 hold2836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 _14406_/X vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2858 _17849_/Q vssd1 vssd1 vccd1 vccd1 hold2858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 _15840_/Q vssd1 vssd1 vccd1 vccd1 hold2869/X sky130_fd_sc_hd__dlygate4sd3_1
X_07875_ _14726_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _18273_/Q hold3835/X _11159_/C vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09545_ hold1994/X _13182_/A _10007_/C vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ hold5910/X _09477_/C _09477_/A vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08427_ _14946_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_403_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08358_ hold944/X _15811_/Q hold134/X vssd1 vssd1 vccd1 vccd1 hold950/A sky130_fd_sc_hd__mux2_1
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08289_ _15513_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _10476_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5440 _11023_/X vssd1 vssd1 vccd1 vccd1 _16831_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10251_ _10830_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5451 _16793_/Q vssd1 vssd1 vccd1 vccd1 hold5451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5462 _11875_/X vssd1 vssd1 vccd1 vccd1 _17115_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5473 _17174_/Q vssd1 vssd1 vccd1 vccd1 hold5473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5484 _10657_/X vssd1 vssd1 vccd1 vccd1 _16709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4750 _09865_/X vssd1 vssd1 vccd1 vccd1 _16445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5495 _16950_/Q vssd1 vssd1 vccd1 vccd1 hold5495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4761 _16445_/Q vssd1 vssd1 vccd1 vccd1 hold4761/X sky130_fd_sc_hd__dlygate4sd3_1
X_10182_ _10560_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10182_/X sky130_fd_sc_hd__or2_1
Xhold4772 _10990_/X vssd1 vssd1 vccd1 vccd1 _16820_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4783 _16417_/Q vssd1 vssd1 vccd1 vccd1 hold4783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4794 _11757_/Y vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14990_ _15205_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout250 _12288_/A vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__buf_4
XFILLER_0_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout261 _11139_/A vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__clkbuf_4
Xfanout272 _13776_/A vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__buf_4
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _17776_/D sky130_fd_sc_hd__and2_1
Xfanout283 _12243_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout294 _12051_/A vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_23_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_23_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16660_ _18216_/CLK _16660_/D vssd1 vssd1 vccd1 vccd1 _16660_/Q sky130_fd_sc_hd__dfxtp_1
X_13872_ hold3791/X _12267_/A _13871_/X vssd1 vssd1 vccd1 vccd1 _13872_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_213_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15611_ _18428_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12823_ hold2579/X hold3179/X _12826_/S vssd1 vssd1 vccd1 vccd1 _12823_/X sky130_fd_sc_hd__mux2_1
X_16591_ _18153_/CLK _16591_/D vssd1 vssd1 vccd1 vccd1 _16591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18330_ _18362_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ hold2188/X _15547_/B _15541_/Y _15548_/C1 vssd1 vssd1 vccd1 vccd1 _15542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12754_ hold1311/X _17429_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__mux2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18293_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ hold2618/X hold4431/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__mux2_1
X_15473_ _15473_/A _15473_/B vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__and2_1
X_12685_ hold1807/X hold4139/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18421_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17212_ _17244_/CLK _17212_/D vssd1 vssd1 vccd1 vccd1 _17212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14424_ hold3069/X _14433_/B _14423_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _14424_/X
+ sky130_fd_sc_hd__o211a_1
X_11636_ hold864/X _17036_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__mux2_1
X_18192_ _18224_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17143_ _17207_/CLK _17143_/D vssd1 vssd1 vccd1 vccd1 _17143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11567_ hold1821/X hold5575/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__mux2_1
X_14355_ _15523_/A hold1476/X hold333/X vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10518_ _10536_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__or2_1
X_13306_ _17589_/Q _17123_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__mux2_1
Xhold709 hold709/A vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17074_ _17889_/CLK _17074_/D vssd1 vssd1 vccd1 vccd1 _17074_/Q sky130_fd_sc_hd__dfxtp_1
X_14286_ hold754/X _14502_/B vssd1 vssd1 vccd1 vccd1 hold755/A sky130_fd_sc_hd__nor2_1
X_11498_ hold1708/X hold4421/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _18411_/CLK _16025_/D vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
X_13237_ _13236_/X hold3555/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10449_ _10998_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ _13161_/X _13167_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17539_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_6_62_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_62_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_12119_ hold2256/X hold4205/X _13862_/C vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17976_ _18040_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
X_13099_ _13098_/X _16905_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux2_1
Xhold1409 _13963_/X vssd1 vssd1 vccd1 vccd1 _17786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16927_ _17808_/CLK _16927_/D vssd1 vssd1 vccd1 vccd1 _16927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16858_ _18032_/CLK _16858_/D vssd1 vssd1 vccd1 vccd1 _16858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15809_ _17426_/CLK _15809_/D vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16789_ _18054_/CLK _16789_/D vssd1 vssd1 vccd1 vccd1 _16789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ hold1603/X _09338_/A2 _09329_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09261_ _15537_/A hold2663/X _09273_/S vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18459_ _18459_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_150_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ hold1910/X _08213_/B _08211_/Y _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08212_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09192_ _15521_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08143_ _08143_/A hold368/X vssd1 vssd1 vccd1 vccd1 hold369/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08074_ _15533_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4002 _16640_/Q vssd1 vssd1 vccd1 vccd1 hold4002/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4013 _13866_/Y vssd1 vssd1 vccd1 vccd1 _13867_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4024 _16356_/Q vssd1 vssd1 vccd1 vccd1 hold4024/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4035 _09811_/X vssd1 vssd1 vccd1 vccd1 _16427_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3301 _17472_/Q vssd1 vssd1 vccd1 vccd1 hold3301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4046 _17067_/Q vssd1 vssd1 vccd1 vccd1 hold4046/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4057 _16885_/Q vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3312 _17585_/Q vssd1 vssd1 vccd1 vccd1 hold3312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4068 _10174_/X vssd1 vssd1 vccd1 vccd1 _16548_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3323 _17385_/Q vssd1 vssd1 vccd1 vccd1 hold3323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3334 _17402_/Q vssd1 vssd1 vccd1 vccd1 hold3334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4079 _17130_/Q vssd1 vssd1 vccd1 vccd1 hold4079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3345 _16473_/Q vssd1 vssd1 vccd1 vccd1 hold3345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2600 _08495_/X vssd1 vssd1 vccd1 vccd1 _15876_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2611 _15805_/Q vssd1 vssd1 vccd1 vccd1 hold2611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3356 _12836_/X vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__buf_6
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2622 _16260_/Q vssd1 vssd1 vccd1 vccd1 hold2622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3367 _17454_/Q vssd1 vssd1 vccd1 vccd1 hold3367/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _12430_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _16105_/D sky130_fd_sc_hd__and2_1
XFILLER_0_215_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2633 _15554_/X vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3378 _12896_/X vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2644 _08457_/X vssd1 vssd1 vccd1 vccd1 _15857_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3389 _09703_/X vssd1 vssd1 vccd1 vccd1 _16391_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1910 _15742_/Q vssd1 vssd1 vccd1 vccd1 hold1910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__buf_4
Xhold2655 _15013_/X vssd1 vssd1 vccd1 vccd1 _18290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 _18172_/Q vssd1 vssd1 vccd1 vccd1 hold1921/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07927_ hold2130/X _07924_/B _07926_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _07927_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2666 _09205_/X vssd1 vssd1 vccd1 vccd1 _16214_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1932 _14763_/X vssd1 vssd1 vccd1 vccd1 _18170_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2677 _16205_/Q vssd1 vssd1 vccd1 vccd1 hold2677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 _14667_/X vssd1 vssd1 vccd1 vccd1 _18124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _18281_/Q vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _18123_/Q vssd1 vssd1 vccd1 vccd1 hold1954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 _15831_/Q vssd1 vssd1 vccd1 vccd1 hold2699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _14697_/X vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ hold1367/X _07869_/B _07857_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _07858_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1976 _14073_/X vssd1 vssd1 vccd1 vccd1 _17839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 _18430_/Q vssd1 vssd1 vccd1 vccd1 hold1987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1998 _17996_/Q vssd1 vssd1 vccd1 vccd1 hold1998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07789_ _07789_/A vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__inv_2
XFILLER_0_196_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _09984_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09463_/C _09463_/D _09458_/Y vssd1 vssd1 vccd1 vccd1 _16313_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12470_ _17328_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11421_ _11652_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14140_ _15213_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14140_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _11553_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11352_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ hold3817/X _10477_/A2 _10302_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14071_ hold1589/X _14107_/A2 _14070_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _11667_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _09494_/A hold957/A _11203_/A vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__a21oi_1
Xhold5270 _17038_/Q vssd1 vssd1 vccd1 vccd1 hold5270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5281 _09886_/X vssd1 vssd1 vccd1 vccd1 _16452_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10234_ hold5082/X _11095_/A2 _10233_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10234_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5292 _17005_/Q vssd1 vssd1 vccd1 vccd1 hold5292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4580 _11962_/X vssd1 vssd1 vccd1 vccd1 _17144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17830_ _17862_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4591 _16008_/Q vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10165_ hold3892/X _10646_/B _10164_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3890 _17559_/Q vssd1 vssd1 vccd1 vccd1 hold3890/X sky130_fd_sc_hd__dlygate4sd3_1
X_17761_ _17890_/CLK _17761_/D vssd1 vssd1 vccd1 vccd1 _17761_/Q sky130_fd_sc_hd__dfxtp_1
X_14973_ hold1638/X _15004_/B _14972_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _14973_/X
+ sky130_fd_sc_hd__o211a_1
X_10096_ hold5711/X _10070_/B _10095_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _10096_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ _18038_/CLK _16712_/D vssd1 vssd1 vccd1 vccd1 _16712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13924_ _15213_/A _17768_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 _13924_/X sky130_fd_sc_hd__mux2_1
X_17692_ _17724_/CLK _17692_/D vssd1 vssd1 vccd1 vccd1 _17692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_396_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17900_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16643_ _18199_/CLK _16643_/D vssd1 vssd1 vccd1 vccd1 _16643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13855_ _13888_/A _13855_/B vssd1 vssd1 vccd1 vccd1 _17738_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_325_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17775_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12806_ hold3333/X _12805_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_186_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16574_ _18220_/CLK _16574_/D vssd1 vssd1 vccd1 vccd1 _16574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10998_ _10998_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _10998_/X sky130_fd_sc_hd__or2_1
X_13786_ hold4461/X _13880_/B _13785_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13786_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18313_ _18319_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 hold844/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15525_ _15525_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ hold3211/X _12736_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12738_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_169_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18276_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15456_ hold854/X _09365_/B _09392_/B hold811/X vssd1 vssd1 vccd1 vccd1 _15456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ hold3770/X _12667_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14910_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18175_ _18175_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _12213_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__or2_1
X_15387_ hold541/X _09357_/A _09386_/D _15896_/Q _15386_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ hold3227/X _12598_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12599_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ _17719_/CLK _17126_/D vssd1 vssd1 vccd1 vccd1 _17126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14338_ _15233_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__or2_1
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold528 la_data_in[30] vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 hold539/A vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17057_ _17871_/CLK _17057_/D vssd1 vssd1 vccd1 vccd1 _17057_/Q sky130_fd_sc_hd__dfxtp_1
X_14269_ hold2265/X _14272_/B _14268_/Y _14538_/C1 vssd1 vssd1 vccd1 vccd1 _14269_/X
+ sky130_fd_sc_hd__o211a_1
X_16008_ _18413_/CLK _16008_/D vssd1 vssd1 vccd1 vccd1 _16008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17129_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08830_ hold454/X hold862/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__mux2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _15852_/Q vssd1 vssd1 vccd1 vccd1 hold1206/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ hold346/X hold727/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold728/A sky130_fd_sc_hd__mux2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _09207_/X vssd1 vssd1 vccd1 vccd1 _16215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17959_ _18059_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _09129_/X vssd1 vssd1 vccd1 vccd1 _16177_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1239 _15582_/Q vssd1 vssd1 vccd1 vccd1 hold1239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08692_ _12386_/A hold538/X vssd1 vssd1 vccd1 vccd1 _15967_/D sky130_fd_sc_hd__and2_1
XFILLER_0_240_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09313_ _15535_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _12768_/A _09244_/B vssd1 vssd1 vccd1 vccd1 _16233_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ hold1587/X _09177_/A2 _09174_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ _14758_/A hold2552/X hold240/X vssd1 vssd1 vccd1 vccd1 _08127_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08057_ hold2601/X _08097_/A2 _08056_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _08057_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3120 _18054_/Q vssd1 vssd1 vccd1 vccd1 hold3120/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3131 _14743_/X vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3142 _14699_/X vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3153 _17350_/Q vssd1 vssd1 vccd1 vccd1 hold3153/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3164 _07798_/X vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3175 _17371_/Q vssd1 vssd1 vccd1 vccd1 hold3175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2430 _17802_/Q vssd1 vssd1 vccd1 vccd1 hold2430/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3186 _14241_/X vssd1 vssd1 vccd1 vccd1 _17919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2441 _15605_/Q vssd1 vssd1 vccd1 vccd1 hold2441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _08322_/X vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3197 _17420_/Q vssd1 vssd1 vccd1 vccd1 hold3197/X sky130_fd_sc_hd__dlygate4sd3_1
X_08959_ hold271/X hold355/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2463 _17868_/Q vssd1 vssd1 vccd1 vccd1 hold2463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 _07917_/X vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1740 _14893_/X vssd1 vssd1 vccd1 vccd1 _18233_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2485 _14597_/X vssd1 vssd1 vccd1 vccd1 _18090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1751 _13890_/X vssd1 vssd1 vccd1 vccd1 _17750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2496 _17927_/Q vssd1 vssd1 vccd1 vccd1 hold2496/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1762 _08000_/X vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11970_ _13794_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__or2_1
Xhold1773 _18222_/Q vssd1 vssd1 vccd1 vccd1 hold1773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _14007_/X vssd1 vssd1 vccd1 vccd1 _17807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1795 _16295_/Q vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10921_ hold4425/X _11207_/B _10920_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10921_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13640_ hold1559/X _17667_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__mux2_1
X_10852_ hold4223/X _11150_/B _10851_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ hold1495/X hold4569/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ hold5108/X _11168_/B _10782_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15310_ hold679/X _09367_/A _09357_/B hold889/X vssd1 vssd1 vccd1 vccd1 _15310_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12531_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _17350_/D sky130_fd_sc_hd__and2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16312_/CLK _16290_/D vssd1 vssd1 vccd1 vccd1 _16290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _09404_/B _15477_/A2 _15487_/B1 hold411/X _15240_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_240_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ hold113/X _12509_/A2 _12507_/A3 _12452_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o311a_1
XFILLER_0_227_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11404_ hold4421/X _12329_/B _11403_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__o211a_1
X_12384_ _12416_/A hold341/X vssd1 vssd1 vccd1 vccd1 _17285_/D sky130_fd_sc_hd__and2_1
X_15172_ hold5976/X _15167_/B hold502/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 hold503/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14123_ hold2240/X _14142_/B _14122_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _14123_/X
+ sky130_fd_sc_hd__o211a_1
X_11335_ hold5018/X _12299_/B _11334_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ hold3934/X _12317_/B _11265_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o211a_1
X_14054_ _14735_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10217_ hold3051/X hold3712/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__mux2_1
X_13005_ _14968_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__or2_1
XTAP_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11197_ _12340_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _16889_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ _18427_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10148_ hold2252/X hold3551/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__mux2_1
XTAP_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _17744_/CLK _17744_/D vssd1 vssd1 vccd1 vccd1 _17744_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ _18073_/Q _16517_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__mux2_1
X_14956_ _15225_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13907_ _13929_/A _13907_/B vssd1 vssd1 vccd1 vccd1 _17759_/D sky130_fd_sc_hd__and2_1
X_17675_ _17707_/CLK _17675_/D vssd1 vssd1 vccd1 vccd1 _17675_/Q sky130_fd_sc_hd__dfxtp_1
X_14887_ hold1519/X _14882_/B _14886_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16626_ _18182_/CLK _16626_/D vssd1 vssd1 vccd1 vccd1 _16626_/Q sky130_fd_sc_hd__dfxtp_1
X_13838_ _13838_/A _13856_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__and3_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16557_ _18113_/CLK _16557_/D vssd1 vssd1 vccd1 vccd1 _16557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13769_ hold2731/X hold4525/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ hold754/X hold533/X vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__or2_4
X_16488_ _18367_/CLK _16488_/D vssd1 vssd1 vccd1 vccd1 _16488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18227_ _18227_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
X_15439_ hold785/X _09386_/A _15437_/X vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18158_ _18216_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17109_ _17153_/CLK _17109_/D vssd1 vssd1 vccd1 vccd1 _17109_/Q sky130_fd_sc_hd__dfxtp_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ _18193_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold336 hold336/A vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold358 data_in[11] vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09931_ hold3203/X _10025_/B _09930_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold369 hold369/A vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout805 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _15007_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout816 _15158_/C1 vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09862_ hold3819/X _10010_/B _09861_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09862_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout827 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14851_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout838 _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/C1 sky130_fd_sc_hd__buf_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _15215_/A vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__buf_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _15414_/A _08813_/B vssd1 vssd1 vccd1 vccd1 _16025_/D sky130_fd_sc_hd__and2_1
Xhold1003 _17946_/Q vssd1 vssd1 vccd1 vccd1 hold1003/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ hold3368/X _10025_/B _09792_/X _14915_/C1 vssd1 vssd1 vccd1 vccd1 _09793_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 input41/X vssd1 vssd1 vccd1 vccd1 hold382/A sky130_fd_sc_hd__buf_1
XFILLER_0_77_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1025 _13029_/X vssd1 vssd1 vccd1 vccd1 _13031_/C sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_247_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18180_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1036 _14980_/X vssd1 vssd1 vccd1 vccd1 hold1036/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1047 input39/X vssd1 vssd1 vccd1 vccd1 hold1047/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _15491_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _15992_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1058 _09137_/X vssd1 vssd1 vccd1 vccd1 _16181_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1069 _14440_/X vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ hold17/X hold265/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08676_/B sky130_fd_sc_hd__mux2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09227_ hold2789/X _09216_/B _09226_/X _12912_/A vssd1 vssd1 vccd1 vccd1 _09227_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ _15541_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_161_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _08137_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ hold2797/X _09106_/B _09088_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _09089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ hold2810/X _16864_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold870 hold870/A vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold881 hold881/A vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 hold892/A vssd1 vssd1 vccd1 vccd1 hold892/X sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ hold1640/X hold4299/X _11147_/C vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _13118_/A _09984_/A _10001_/X vssd1 vssd1 vccd1 vccd1 _10002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2260 _18161_/Q vssd1 vssd1 vccd1 vccd1 hold2260/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _14988_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__or2_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2271 _17851_/Q vssd1 vssd1 vccd1 vccd1 hold2271/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2282 _15662_/Q vssd1 vssd1 vccd1 vccd1 hold2282/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _17658_/CLK _15790_/D vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2293 _17837_/Q vssd1 vssd1 vccd1 vccd1 hold2293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1570 _14725_/X vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14741_ hold1962/X _14774_/B _14740_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14741_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 _18255_/Q vssd1 vssd1 vccd1 vccd1 hold1581/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1592 _14917_/X vssd1 vssd1 vccd1 vccd1 _18243_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ hold3506/X _12374_/B _11952_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _11953_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10904_ hold2647/X _16792_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10905_/B sky130_fd_sc_hd__mux2_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17482_/CLK _17460_/D vssd1 vssd1 vccd1 vccd1 _17460_/Q sky130_fd_sc_hd__dfxtp_1
X_14672_ _14726_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__or2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ hold4173/X _13871_/B _11883_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _18322_/CLK _16411_/D vssd1 vssd1 vccd1 vccd1 _16411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13623_ _13623_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17391_ _18455_/CLK _17391_/D vssd1 vssd1 vccd1 vccd1 _17391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10835_ hold1741/X _16769_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16342_ _18393_/CLK _16342_/D vssd1 vssd1 vccd1 vccd1 _16342_/Q sky130_fd_sc_hd__dfxtp_1
X_13554_ _13746_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ _17947_/Q _16746_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__mux2_1
X_12505_ hold20/X _08597_/Y _08868_/X _12504_/X _09063_/A vssd1 vssd1 vccd1 vccd1
+ hold21/A sky130_fd_sc_hd__o311a_1
XFILLER_0_164_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16273_ _17517_/CLK _16273_/D vssd1 vssd1 vccd1 vccd1 _16273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ hold3128/X hold4664/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__mux2_1
X_13485_ _13776_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _18012_/CLK hold912/X vssd1 vssd1 vccd1 vccd1 hold911/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ hold5988/X _15219_/B hold973/X _15024_/A vssd1 vssd1 vccd1 vccd1 hold974/A
+ sky130_fd_sc_hd__o211a_1
X_12436_ _12436_/A hold146/X vssd1 vssd1 vccd1 vccd1 _17311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15155_ _15209_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12367_ _12367_/A _12367_/B vssd1 vssd1 vccd1 vccd1 _17279_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ _15233_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ hold2314/X _16930_/Q _11480_/S vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15086_ hold2746/X _15113_/B _15085_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ _13825_/A _12298_/B vssd1 vssd1 vccd1 vccd1 _17256_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_240_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ hold2031/X _14038_/B _14036_/Y _14376_/A vssd1 vssd1 vccd1 vccd1 _14037_/X
+ sky130_fd_sc_hd__o211a_1
X_11249_ hold1752/X hold3600/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_340_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17283_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15988_ _18300_/CLK _15988_/D vssd1 vssd1 vccd1 vccd1 hold440/A sky130_fd_sc_hd__dfxtp_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17727_ _17729_/CLK _17727_/D vssd1 vssd1 vccd1 vccd1 _17727_/Q sky130_fd_sc_hd__dfxtp_1
X_14939_ hold1599/X _14946_/B _14938_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _14854_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17658_ _17658_/CLK _17658_/D vssd1 vssd1 vccd1 vccd1 _17658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16609_ _18229_/CLK _16609_/D vssd1 vssd1 vccd1 vccd1 _16609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08391_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _15827_/D sky130_fd_sc_hd__and2_1
XFILLER_0_212_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17589_ _17650_/CLK _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ hold47/X hold417/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5803 hold5940/X vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 hold309/X vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5814 output95/X vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_12
XFILLER_0_182_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5825 output96/X vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5836 hold5836/A vssd1 vssd1 vccd1 vccd1 hold5836/X sky130_fd_sc_hd__buf_2
Xhold5847 _18412_/Q vssd1 vssd1 vccd1 vccd1 hold5847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__clkbuf_2
Xhold133 hold204/X vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5858 hold5858/A vssd1 vssd1 vccd1 vccd1 hold5858/X sky130_fd_sc_hd__clkbuf_4
Xhold144 input24/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__buf_1
XFILLER_0_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5869 _18410_/Q vssd1 vssd1 vccd1 vccd1 hold5869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_428_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09914_ hold1387/X _16462_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__mux2_1
Xfanout602 _09366_/Y vssd1 vssd1 vccd1 vccd1 _15484_/B1 sky130_fd_sc_hd__buf_6
Xhold199 hold528/X vssd1 vssd1 vccd1 vccd1 hold529/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 _09358_/Y vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__clkbuf_8
Xfanout624 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15490_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout635 hold5897/X vssd1 vssd1 vccd1 vccd1 _13304_/B1 sky130_fd_sc_hd__buf_8
XFILLER_0_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout646 _13714_/C1 vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__buf_2
X_09845_ hold2238/X hold3672/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__mux2_1
Xfanout657 _12987_/A vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__clkbuf_2
Xfanout668 _13801_/C1 vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__buf_4
Xfanout679 fanout692/X vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__buf_2
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09776_ hold1646/X _16416_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ hold150/X _15985_/Q _08727_/S vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _12404_/A hold873/X vssd1 vssd1 vccd1 vccd1 _15951_/D sky130_fd_sc_hd__and2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _12408_/A hold336/X vssd1 vssd1 vccd1 vccd1 _15918_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ hold4701/X _10524_/A _10619_/X vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10551_ _10998_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__or2_1
X_13270_ _13270_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ hold2880/X _17231_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _12222_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ hold1456/X _17208_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18337_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11103_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12083_ hold3102/X hold4401/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__mux2_1
X_16960_ _17891_/CLK _16960_/D vssd1 vssd1 vccd1 vccd1 _16960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _16089_/CLK _15911_/D vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__dfxtp_1
X_11034_ _11121_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__or2_1
X_16891_ _18060_/CLK _16891_/D vssd1 vssd1 vccd1 vccd1 _16891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _17739_/CLK _15842_/D vssd1 vssd1 vccd1 vccd1 _15842_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _16180_/Q vssd1 vssd1 vccd1 vccd1 hold2090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _17724_/CLK _15773_/D vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12985_ hold2102/X _17506_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__mux2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _18398_/CLK _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _15225_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__or2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ hold2267/X hold5360/X _13793_/S vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__mux2_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17443_ _17444_/CLK _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14655_ hold1927/X _14666_/B _14654_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14655_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11867_ hold2438/X hold3596/X _13868_/C vssd1 vssd1 vccd1 vccd1 _11868_/B sky130_fd_sc_hd__mux2_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13606_ hold4225/X _13802_/B _13605_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__o211a_1
X_17374_ _17376_/CLK _17374_/D vssd1 vssd1 vccd1 vccd1 _17374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ _11106_/A _10818_/B vssd1 vssd1 vccd1 vccd1 _10818_/X sky130_fd_sc_hd__or2_1
X_14586_ _14910_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _17090_/Q _12344_/B _12344_/C vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16325_ _18300_/CLK _16325_/D vssd1 vssd1 vccd1 vccd1 _16325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13537_ hold5747/X _13832_/B _13536_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10749_ _11064_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16256_ _17378_/CLK _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Q sky130_fd_sc_hd__dfxtp_1
X_13468_ hold4243/X _13883_/B _13467_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15207_ _15207_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__or2_1
X_12419_ hold402/X hold830/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold831/A sky130_fd_sc_hd__mux2_1
XFILLER_0_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16187_ _17506_/CLK _16187_/D vssd1 vssd1 vccd1 vccd1 _16187_/Q sky130_fd_sc_hd__dfxtp_1
X_13399_ hold4483/X _13877_/B _13398_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _13399_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4409 _17143_/Q vssd1 vssd1 vccd1 vccd1 hold4409/X sky130_fd_sc_hd__dlygate4sd3_1
X_15138_ hold2238/X _15167_/B _15137_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3708 _16385_/Q vssd1 vssd1 vccd1 vccd1 hold3708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3719 _10246_/X vssd1 vssd1 vccd1 vccd1 _16572_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15069_ hold719/A _18318_/Q _15069_/S vssd1 vssd1 vccd1 vccd1 hold623/A sky130_fd_sc_hd__mux2_1
X_07960_ _15529_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07960_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07891_ hold1373/X _07918_/B _07890_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07891_/X
+ sky130_fd_sc_hd__o211a_1
X_09630_ _09933_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09561_ _11097_/A _09561_/B vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08512_ hold2500/X _08503_/Y _08511_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08512_/X
+ sky130_fd_sc_hd__o211a_1
X_09492_ _13029_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _09494_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ _14443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08374_ hold246/A _15819_/Q hold134/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5600 _12052_/X vssd1 vssd1 vccd1 vccd1 _17174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5611 _16826_/Q vssd1 vssd1 vccd1 vccd1 hold5611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5622 _09640_/X vssd1 vssd1 vccd1 vccd1 _16370_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5633 _16769_/Q vssd1 vssd1 vccd1 vccd1 hold5633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5644 _11032_/X vssd1 vssd1 vccd1 vccd1 _16834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4910 _10222_/X vssd1 vssd1 vccd1 vccd1 _16564_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5655 _16350_/Q vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4921 _16573_/Q vssd1 vssd1 vccd1 vccd1 hold4921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5666 _10192_/X vssd1 vssd1 vccd1 vccd1 _16554_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4932 _16693_/Q vssd1 vssd1 vccd1 vccd1 hold4932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5677 _16446_/Q vssd1 vssd1 vccd1 vccd1 hold5677/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4943 _10519_/X vssd1 vssd1 vccd1 vccd1 _16663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5688 _10078_/X vssd1 vssd1 vccd1 vccd1 _16516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_262_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17960_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_218_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4954 _16661_/Q vssd1 vssd1 vccd1 vccd1 hold4954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5699 _16514_/Q vssd1 vssd1 vccd1 vccd1 hold5699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4965 _12286_/X vssd1 vssd1 vccd1 vccd1 _17252_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4976 _17128_/Q vssd1 vssd1 vccd1 vccd1 hold4976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4987 _10447_/X vssd1 vssd1 vccd1 vccd1 _16639_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout410 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__buf_6
Xfanout421 _13996_/B vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__clkbuf_8
Xfanout432 _13622_/S vssd1 vssd1 vccd1 vccd1 _13808_/C sky130_fd_sc_hd__clkbuf_8
Xhold4998 _16927_/Q vssd1 vssd1 vccd1 vccd1 hold4998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout443 _13622_/S vssd1 vssd1 vccd1 vccd1 _12029_/S sky130_fd_sc_hd__clkbuf_4
Xfanout454 _11168_/C vssd1 vssd1 vccd1 vccd1 _11738_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout465 _13874_/C vssd1 vssd1 vccd1 vccd1 _13886_/C sky130_fd_sc_hd__buf_6
Xfanout476 _11480_/S vssd1 vssd1 vccd1 vccd1 _12344_/C sky130_fd_sc_hd__clkbuf_8
X_09828_ _09933_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__or2_1
Xfanout487 _11057_/S vssd1 vssd1 vccd1 vccd1 _09824_/S sky130_fd_sc_hd__clkbuf_4
Xfanout498 _11096_/S vssd1 vssd1 vccd1 vccd1 _10580_/C sky130_fd_sc_hd__buf_6
Xclkbuf_6_13_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_13_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ _09954_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__or2_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ hold3750/X _12769_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ hold4679/X _12204_/A _11720_/X vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ hold5990/X _14433_/B hold1068/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14440_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _16691_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ _15105_/A hold2545/X hold333/X vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__mux2_1
X_11583_ _11679_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16110_ _17523_/CLK _16110_/D vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13322_ hold2500/X _17561_/Q _13622_/S vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10534_ hold4867/X _10628_/B _10533_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10534_/X
+ sky130_fd_sc_hd__o211a_1
X_17090_ _17904_/CLK _17090_/D vssd1 vssd1 vccd1 vccd1 _17090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _17297_/CLK _16041_/D vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ hold5070/X _10565_/B _10464_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__o211a_1
X_13253_ _13252_/X hold3551/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__or2_1
X_13184_ _13177_/X _13183_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17541_/D sky130_fd_sc_hd__o21a_1
X_10396_ hold5240/X _10625_/B _10395_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_52_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_52_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_206_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12135_ _12267_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__or2_1
X_17992_ _18230_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16943_ _17821_/CLK _16943_/D vssd1 vssd1 vccd1 vccd1 _16943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _13794_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ hold4467/X _11768_/B _11016_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__o211a_1
X_16874_ _18430_/CLK _16874_/D vssd1 vssd1 vccd1 vccd1 _16874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ _17738_/CLK _15825_/D vssd1 vssd1 vccd1 vccd1 _15825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ _17702_/CLK _15756_/D vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ hold3171/X _12967_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18459_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ hold3006/X _14714_/B _14706_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14707_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11919_ _13716_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15687_ _17179_/CLK _15687_/D vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ hold3394/X _12898_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__mux2_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17426_ _17426_/CLK _17426_/D vssd1 vssd1 vccd1 vccd1 _17426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _15193_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17357_ _17378_/CLK _17357_/D vssd1 vssd1 vccd1 vccd1 _17357_/Q sky130_fd_sc_hd__dfxtp_1
X_14569_ _15193_/A _14557_/Y hold2110/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16308_ _16312_/CLK _16308_/D vssd1 vssd1 vccd1 vccd1 _16308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _15549_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08090_/X sky130_fd_sc_hd__or2_1
X_17288_ _17301_/CLK _17288_/D vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16239_ _17420_/CLK _16239_/D vssd1 vssd1 vccd1 vccd1 _16239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4206 _12025_/X vssd1 vssd1 vccd1 vccd1 _17165_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4217 _17202_/Q vssd1 vssd1 vccd1 vccd1 hold4217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4228 _11539_/X vssd1 vssd1 vccd1 vccd1 _17003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4239 _10672_/X vssd1 vssd1 vccd1 vccd1 _16714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3505 _13375_/X vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3516 _10771_/X vssd1 vssd1 vccd1 vccd1 _16747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3527 _17391_/Q vssd1 vssd1 vccd1 vccd1 hold3527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08992_ _12430_/A hold170/X vssd1 vssd1 vccd1 vccd1 _16113_/D sky130_fd_sc_hd__and2_1
Xhold3538 _10044_/Y vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3549 _16535_/Q vssd1 vssd1 vccd1 vccd1 hold3549/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_76_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2804 _17801_/Q vssd1 vssd1 vccd1 vccd1 hold2804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 _14496_/X vssd1 vssd1 vccd1 vccd1 _18043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2826 _18153_/Q vssd1 vssd1 vccd1 vccd1 hold2826/X sky130_fd_sc_hd__dlygate4sd3_1
X_07943_ hold1221/X _07991_/A2 _07942_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _07943_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2837 _08310_/X vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2848 _16179_/Q vssd1 vssd1 vccd1 vccd1 hold2848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2859 _14093_/X vssd1 vssd1 vccd1 vccd1 _17849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07874_ hold1239/X _07869_/B _07873_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ hold3399/X _10013_/B _09612_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09613_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ hold5571/X _09832_/A2 _09543_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09475_ hold5910/X _09477_/C _09474_/Y vssd1 vssd1 vccd1 vccd1 _16319_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08426_ hold5995/X _08433_/B hold1086/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08357_ _12741_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _15810_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08288_ hold1495/X _08336_/A2 _08287_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08288_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_443_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17693_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5430 _10690_/X vssd1 vssd1 vccd1 vccd1 _16720_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10250_ hold2787/X _16574_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5441 _17078_/Q vssd1 vssd1 vccd1 vccd1 hold5441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5452 _10813_/X vssd1 vssd1 vccd1 vccd1 _16761_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5463 _16740_/Q vssd1 vssd1 vccd1 vccd1 hold5463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5474 _11956_/X vssd1 vssd1 vccd1 vccd1 _17142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4740 _09847_/X vssd1 vssd1 vccd1 vccd1 _16439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5485 _16843_/Q vssd1 vssd1 vccd1 vccd1 hold5485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ hold1855/X hold4773/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__mux2_1
Xhold5496 _11284_/X vssd1 vssd1 vccd1 vccd1 _16918_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4751 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold4751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4762 _09769_/X vssd1 vssd1 vccd1 vccd1 _16413_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4773 _16551_/Q vssd1 vssd1 vccd1 vccd1 hold4773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4784 _09685_/X vssd1 vssd1 vccd1 vccd1 _16385_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4795 _16517_/Q vssd1 vssd1 vccd1 vccd1 hold4795/X sky130_fd_sc_hd__buf_2
Xfanout240 _10477_/A2 vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__buf_4
XFILLER_0_206_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout251 _13623_/A vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__clkbuf_4
Xfanout262 _11139_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__buf_4
Xfanout273 fanout334/X vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__clkbuf_4
X_13940_ _14782_/A hold2314/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout284 _12051_/A vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__buf_4
Xfanout295 fanout334/X vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__buf_4
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _17744_/Q _13871_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13871_/X sky130_fd_sc_hd__and3_1
XFILLER_0_202_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15610_ _17258_/CLK _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
X_12822_ _12894_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _17450_/D sky130_fd_sc_hd__and2_1
X_16590_ _18178_/CLK _16590_/D vssd1 vssd1 vccd1 vccd1 _16590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12753_ _12759_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _17427_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18292_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11704_ hold4515/X _12344_/B _11703_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11704_/X
+ sky130_fd_sc_hd__o211a_1
X_15472_ _15481_/A1 _15465_/X _15471_/X _15481_/B1 hold5888/A vssd1 vssd1 vccd1 vccd1
+ _15472_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_155_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12780_/A _12684_/B vssd1 vssd1 vccd1 vccd1 _17404_/D sky130_fd_sc_hd__and2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17590_/CLK _17211_/D vssd1 vssd1 vccd1 vccd1 _17211_/Q sky130_fd_sc_hd__dfxtp_1
X_14423_ _15103_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14423_/X sky130_fd_sc_hd__or2_1
X_18191_ _18223_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11635_ hold4046/X _11729_/B _11634_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11635_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17142_ _17210_/CLK _17142_/D vssd1 vssd1 vccd1 vccd1 _17142_/Q sky130_fd_sc_hd__dfxtp_1
X_14354_ _14368_/A _14354_/B vssd1 vssd1 vccd1 vccd1 _17974_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11566_ hold5545/X _11762_/B _11565_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_184_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18202_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13305_ _13305_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13305_/X sky130_fd_sc_hd__and2_1
XFILLER_0_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10517_ hold2967/X hold3990/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17073_ _17887_/CLK _17073_/D vssd1 vssd1 vccd1 vccd1 _17073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14285_ hold5992/X _14266_/B hold602/X _14370_/A vssd1 vssd1 vccd1 vccd1 hold603/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ hold5371/X _12329_/B _11496_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11497_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ _17347_/CLK _16024_/D vssd1 vssd1 vccd1 vccd1 _16024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ hold4676/X _13235_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ hold1839/X _16640_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_237_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _13311_/A1 _13165_/X _13166_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13167_/X
+ sky130_fd_sc_hd__o211a_1
X_10379_ hold2852/X _16617_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12118_ hold5150/X _13798_/A2 _12117_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13098_ _17563_/Q _17097_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17975_ _17975_/CLK _17975_/D vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12049_ hold3460/X _12274_/A2 _12048_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12049_/X
+ sky130_fd_sc_hd__o211a_1
X_16926_ _17899_/CLK _16926_/D vssd1 vssd1 vccd1 vccd1 _16926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16857_ _18058_/CLK _16857_/D vssd1 vssd1 vccd1 vccd1 _16857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15808_ _17724_/CLK _15808_/D vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _18053_/CLK _16788_/D vssd1 vssd1 vccd1 vccd1 _16788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ _17742_/CLK _15739_/D vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09260_ _12738_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__and2_1
X_18458_ _18460_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08211_ _15004_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _17431_/CLK _17409_/D vssd1 vssd1 vccd1 vccd1 _17409_/Q sky130_fd_sc_hd__dfxtp_1
X_09191_ hold1050/X _09216_/B _09190_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _09191_/X
+ sky130_fd_sc_hd__o211a_1
X_18389_ _18389_/CLK hold965/X vssd1 vssd1 vccd1 vccd1 hold964/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ hold367/X _15710_/Q hold240/X vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__mux2_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08073_ hold2267/X _08097_/A2 _08072_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _08073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4003 _10354_/X vssd1 vssd1 vccd1 vccd1 _16608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4014 _17065_/Q vssd1 vssd1 vccd1 vccd1 hold4014/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4025 _09502_/X vssd1 vssd1 vccd1 vccd1 _16324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4036 _16433_/Q vssd1 vssd1 vccd1 vccd1 hold4036/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3302 _17443_/Q vssd1 vssd1 vccd1 vccd1 hold3302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4047 _11635_/X vssd1 vssd1 vccd1 vccd1 _17035_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4058 _11089_/X vssd1 vssd1 vccd1 vccd1 _16853_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3313 _13875_/Y vssd1 vssd1 vccd1 vccd1 _13876_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3324 _12626_/X vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4069 _16939_/Q vssd1 vssd1 vccd1 vccd1 hold4069/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3335 _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3346 _09853_/X vssd1 vssd1 vccd1 vccd1 _16441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2601 _15668_/Q vssd1 vssd1 vccd1 vccd1 hold2601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2612 _15684_/Q vssd1 vssd1 vccd1 vccd1 hold2612/X sky130_fd_sc_hd__dlygate4sd3_1
X_08975_ hold353/X hold457/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3357 _16425_/Q vssd1 vssd1 vccd1 vccd1 hold3357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3368 _16453_/Q vssd1 vssd1 vccd1 vccd1 hold3368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 _09300_/X vssd1 vssd1 vccd1 vccd1 _16260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkbuf_2
Xhold3379 _16495_/Q vssd1 vssd1 vccd1 vccd1 hold3379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _18031_/Q vssd1 vssd1 vccd1 vccd1 hold2634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1900 _14579_/X vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2645 _15616_/Q vssd1 vssd1 vccd1 vccd1 hold2645/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1911 _08212_/X vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _15549_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__or2_1
Xhold2656 _15657_/Q vssd1 vssd1 vccd1 vccd1 hold2656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 _14767_/X vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2667 _15601_/Q vssd1 vssd1 vccd1 vccd1 hold2667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__buf_4
Xhold1933 _18209_/Q vssd1 vssd1 vccd1 vccd1 hold1933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 _09187_/X vssd1 vssd1 vccd1 vccd1 _16205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _18137_/Q vssd1 vssd1 vccd1 vccd1 hold2689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1944 _14995_/X vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 _14665_/X vssd1 vssd1 vccd1 vccd1 _18123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1966 _18286_/Q vssd1 vssd1 vccd1 vccd1 hold1966/X sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _14529_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07857_/X sky130_fd_sc_hd__or2_1
Xhold1977 _18217_/Q vssd1 vssd1 vccd1 vccd1 hold1977/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1988 _17960_/Q vssd1 vssd1 vccd1 vccd1 hold1988/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1999 _14400_/X vssd1 vssd1 vccd1 vccd1 _17996_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07788_ _07788_/A vssd1 vssd1 vccd1 vccd1 _07788_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ hold1799/X _16333_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09463_/C _09463_/D _09440_/X vssd1 vssd1 vccd1 vccd1 _09458_/Y sky130_fd_sc_hd__a21boi_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _15523_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08409_/X sky130_fd_sc_hd__or2_1
X_09389_ _07805_/A _09362_/A _09362_/D vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11420_ hold1210/X _16964_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11351_ hold3061/X _16941_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10476_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14070_ _14517_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ hold2233/X hold4815/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__mux2_1
Xhold5260 _16562_/Q vssd1 vssd1 vccd1 vccd1 hold5260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _13048_/A hold920/X hold819/X vssd1 vssd1 vccd1 vccd1 hold956/A sky130_fd_sc_hd__a21o_1
X_10233_ _10830_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5271 _11548_/X vssd1 vssd1 vccd1 vccd1 _17006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5282 _17645_/Q vssd1 vssd1 vccd1 vccd1 hold5282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5293 _11449_/X vssd1 vssd1 vccd1 vccd1 _16973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4570 _13477_/X vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4581 hold5881/X vssd1 vssd1 vccd1 vccd1 hold5882/A sky130_fd_sc_hd__buf_4
X_10164_ _10998_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__or2_1
Xhold4592 _15393_/X vssd1 vssd1 vccd1 vccd1 _15394_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3880 _16371_/Q vssd1 vssd1 vccd1 vccd1 hold3880/X sky130_fd_sc_hd__dlygate4sd3_1
X_14972_ _14972_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or2_1
X_10095_ _10191_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__or2_1
Xhold3891 _13798_/X vssd1 vssd1 vccd1 vccd1 _17719_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17760_ _17889_/CLK _17760_/D vssd1 vssd1 vccd1 vccd1 _17760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16711_ _18012_/CLK _16711_/D vssd1 vssd1 vccd1 vccd1 _16711_/Q sky130_fd_sc_hd__dfxtp_1
X_13923_ _13923_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _17767_/D sky130_fd_sc_hd__and2_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17691_ _17723_/CLK _17691_/D vssd1 vssd1 vccd1 vccd1 _17691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16642_ _18230_/CLK _16642_/D vssd1 vssd1 vccd1 vccd1 _16642_/Q sky130_fd_sc_hd__dfxtp_1
X_13854_ hold3637/X _13779_/A _13853_/X vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12805_ hold2665/X hold3330/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16573_ _18225_/CLK _16573_/D vssd1 vssd1 vccd1 vccd1 _16573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _13791_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13785_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10997_ hold2367/X _16823_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18312_ _18323_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_15524_ hold1237/X _15560_/A2 _15523_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _15524_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ hold2531/X hold3199/X _12748_/S vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_365_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17712_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18243_ _18303_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15455_ _15455_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12667_ hold2518/X _17400_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14406_ hold2846/X _14446_/A2 _14405_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14406_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18174_ _18287_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11618_ hold2278/X hold5088/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__mux2_1
X_15386_ _17342_/Q _15479_/B1 _09362_/D _16119_/Q vssd1 vssd1 vccd1 vccd1 _15386_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12598_ hold1603/X _17377_/Q _12967_/S vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__mux2_1
X_17125_ _17253_/CLK _17125_/D vssd1 vssd1 vccd1 vccd1 _17125_/Q sky130_fd_sc_hd__dfxtp_1
X_14337_ hold1307/X _14326_/B _14336_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14337_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11549_ hold2776/X _17007_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold507 hold507/A vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 hold518/A vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold529 hold529/A vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _17905_/CLK _17056_/D vssd1 vssd1 vccd1 vccd1 _17056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14268_ _14878_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__nand2_1
X_16007_ _18413_/CLK _16007_/D vssd1 vssd1 vccd1 vccd1 hold422/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13219_ _13218_/X _16920_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ hold2197/X _14198_/B _14198_/Y _08117_/A vssd1 vssd1 vccd1 vccd1 _14199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1207 _08444_/X vssd1 vssd1 vccd1 vccd1 _15852_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08760_ _12412_/A hold815/X vssd1 vssd1 vccd1 vccd1 _16000_/D sky130_fd_sc_hd__and2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _18072_/Q vssd1 vssd1 vccd1 vccd1 hold1218/X sky130_fd_sc_hd__dlygate4sd3_1
X_17958_ _18124_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1229 _18206_/Q vssd1 vssd1 vccd1 vccd1 hold1229/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17365_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _17883_/CLK _16909_/D vssd1 vssd1 vccd1 vccd1 _16909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ hold454/X hold537/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold538/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17889_ _17889_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ hold2993/X _09325_/B _09311_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09312_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ _15519_/A hold1121/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09243_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ _15557_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08125_ _08125_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _15701_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08056_ _15515_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3110 _17956_/Q vssd1 vssd1 vccd1 vccd1 hold3110/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3121 _14520_/X vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3132 _18028_/Q vssd1 vssd1 vccd1 vccd1 hold3132/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3143 _18166_/Q vssd1 vssd1 vccd1 vccd1 hold3143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3154 _12521_/X vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3165 _17925_/Q vssd1 vssd1 vccd1 vccd1 hold3165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2420 _15851_/Q vssd1 vssd1 vccd1 vccd1 hold2420/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3176 _12584_/X vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2431 _13995_/X vssd1 vssd1 vccd1 vccd1 _17802_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _12426_/A hold784/X vssd1 vssd1 vccd1 vccd1 _16096_/D sky130_fd_sc_hd__and2_1
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2442 _07923_/X vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3187 _17449_/Q vssd1 vssd1 vccd1 vccd1 hold3187/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2453 _17915_/Q vssd1 vssd1 vccd1 vccd1 hold2453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3198 _12731_/X vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 _14133_/X vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2475 _15882_/Q vssd1 vssd1 vccd1 vccd1 hold2475/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1730 _14131_/X vssd1 vssd1 vccd1 vccd1 _17867_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ hold2422/X _07918_/B _07908_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _07909_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2486 _15661_/Q vssd1 vssd1 vccd1 vccd1 hold2486/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1741 _17970_/Q vssd1 vssd1 vccd1 vccd1 hold1741/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _17753_/Q vssd1 vssd1 vccd1 vccd1 hold1752/X sky130_fd_sc_hd__dlygate4sd3_1
X_08889_ _12408_/A hold315/X vssd1 vssd1 vccd1 vccd1 _16062_/D sky130_fd_sc_hd__and2_1
Xhold2497 _14257_/X vssd1 vssd1 vccd1 vccd1 _17927_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1763 _17871_/Q vssd1 vssd1 vccd1 vccd1 hold1763/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1774 _14871_/X vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1785 _15664_/Q vssd1 vssd1 vccd1 vccd1 hold1785/X sky130_fd_sc_hd__dlygate4sd3_1
X_10920_ _11124_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__or2_1
XFILLER_0_224_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1796 _09419_/X vssd1 vssd1 vccd1 vccd1 _16295_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _11637_/A _10851_/B vssd1 vssd1 vccd1 vccd1 _10851_/X sky130_fd_sc_hd__or2_1
XFILLER_0_212_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ hold4511/X _13847_/B _13569_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13570_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _11643_/A _10782_/B vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__or2_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12521_ hold3153/X _12520_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ hold634/X _15486_/A2 _09357_/B hold661/X vssd1 vssd1 vccd1 vccd1 _15240_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _17319_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11403_ _12234_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__or2_1
X_15171_ hold559/A _15171_/B vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12383_ hold312/X hold340/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold341/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _14246_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14122_/X sky130_fd_sc_hd__or2_1
X_11334_ _12204_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ hold2802/X _14038_/B _14052_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14053_/X
+ sky130_fd_sc_hd__o211a_1
X_11265_ _12285_/A _11265_/B vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5090 _16478_/Q vssd1 vssd1 vccd1 vccd1 hold5090/X sky130_fd_sc_hd__dlygate4sd3_1
X_13004_ _14897_/A hold533/A vssd1 vssd1 vccd1 vccd1 _13017_/B sky130_fd_sc_hd__or2_2
XFILLER_0_24_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10216_ hold4727/X _10598_/B _10215_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10216_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11196_ hold4881/X _11115_/A _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ _17876_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10147_ hold3677/X _10477_/A2 _10146_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14955_ hold984/X _14946_/B _14954_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 hold985/A
+ sky130_fd_sc_hd__o211a_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _17744_/CLK _17743_/D vssd1 vssd1 vccd1 vccd1 _17743_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ hold5687/X _10598_/B _10077_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _10078_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13906_ _14246_/A hold2169/X hold124/X vssd1 vssd1 vccd1 vccd1 _13907_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14886_ _15225_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14886_/X sky130_fd_sc_hd__or2_1
X_17674_ _17740_/CLK _17674_/D vssd1 vssd1 vccd1 vccd1 _17674_/Q sky130_fd_sc_hd__dfxtp_1
X_16625_ _18213_/CLK _16625_/D vssd1 vssd1 vccd1 vccd1 _16625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13837_ _13873_/A _13837_/B vssd1 vssd1 vccd1 vccd1 _17732_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16556_ _18176_/CLK _16556_/D vssd1 vssd1 vccd1 vccd1 _16556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ hold5749/X _13862_/B _13767_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _13768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12719_ hold3693/X _12718_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__mux2_1
X_15507_ hold754/X hold533/X vssd1 vssd1 vccd1 vccd1 _15507_/Y sky130_fd_sc_hd__nor2_4
X_16487_ _18272_/CLK _16487_/D vssd1 vssd1 vccd1 vccd1 _16487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ hold5238/X _13817_/B _13698_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15438_ hold613/X _09367_/A _15479_/B1 _17347_/Q vssd1 vssd1 vccd1 vccd1 _15438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18226_ _18226_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18157_ _18163_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
X_15369_ hold633/X _15485_/A2 _15488_/A2 hold493/X _15368_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17108_ _17711_/CLK _17108_/D vssd1 vssd1 vccd1 vccd1 _17108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold315 hold315/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _18224_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold337 hold337/A vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09930_ _11061_/A _09930_/B vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__or2_1
X_17039_ _17834_/CLK _17039_/D vssd1 vssd1 vccd1 vccd1 _17039_/Q sky130_fd_sc_hd__dfxtp_1
Xhold359 hold22/X vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout806 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout817 _15026_/A vssd1 vssd1 vccd1 vccd1 _15158_/C1 sky130_fd_sc_hd__clkbuf_8
X_09861_ _09933_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__buf_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout839 _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14869_/C1 sky130_fd_sc_hd__buf_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ hold88/X hold91/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09984_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__or2_1
Xhold1004 _14297_/X vssd1 vssd1 vccd1 vccd1 _17946_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 hold382/X vssd1 vssd1 vccd1 vccd1 hold1015/X sky130_fd_sc_hd__buf_4
Xhold1026 _16150_/Q vssd1 vssd1 vccd1 vccd1 hold1026/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1037 _14981_/X vssd1 vssd1 vccd1 vccd1 _18274_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ hold47/X hold722/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__mux2_1
Xhold1048 _15151_/X vssd1 vssd1 vccd1 vccd1 hold1048/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1059 _15807_/Q vssd1 vssd1 vccd1 vccd1 hold1059/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _09015_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _15958_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_287_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17996_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_216_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _15555_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ hold2739/X _09164_/B _09156_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08108_ _15513_/A hold2671/X hold240/X vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _14988_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _14726_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08039_/X sky130_fd_sc_hd__or2_1
Xhold860 hold860/A vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 hold871/A vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold882 hold882/A vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 hold893/A vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ hold4415/X _11147_/B _11049_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _11050_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10001_ _16491_/Q _10025_/B _10001_/C vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 _18376_/Q vssd1 vssd1 vccd1 vccd1 hold2250/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2261 _14745_/X vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2272 _14097_/X vssd1 vssd1 vccd1 vccd1 _17851_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2283 _08042_/X vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _14069_/X vssd1 vssd1 vccd1 vccd1 _17837_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _08334_/X vssd1 vssd1 vccd1 vccd1 _15800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 _18356_/Q vssd1 vssd1 vccd1 vccd1 hold1571/X sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ _14794_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _12273_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1582 _14941_/X vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1593 _17916_/Q vssd1 vssd1 vccd1 vccd1 hold1593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10903_ hold3922/X _10646_/B _10902_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10903_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14671_ hold1513/X _14666_/B _14670_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14671_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _12267_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _18353_/CLK _16410_/D vssd1 vssd1 vccd1 vccd1 _16410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ hold2451/X _17661_/Q _13622_/S vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__mux2_1
X_10834_ hold5204/X _11216_/B _10833_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10834_/X
+ sky130_fd_sc_hd__o211a_1
X_17390_ _18455_/CLK _17390_/D vssd1 vssd1 vccd1 vccd1 _17390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _18356_/CLK _16341_/D vssd1 vssd1 vccd1 vccd1 _16341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13553_ hold1006/X hold4348/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__mux2_1
X_10765_ hold4385/X _11147_/B _10764_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10765_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _17345_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16272_ _17376_/CLK hold906/X vssd1 vssd1 vccd1 vccd1 hold905/A sky130_fd_sc_hd__dfxtp_1
X_13484_ hold1206/X _17615_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__mux2_1
X_10696_ hold4295/X _11753_/B _10695_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15223_ hold972/X _15233_/B vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__or2_1
X_18011_ _18043_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
X_12435_ hold145/X _17311_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__mux2_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ hold1466/X _15165_/B _15153_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ hold3734/X _12246_/A _12365_/X vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14105_ hold1620/X _14107_/A2 _14104_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _14105_/X
+ sky130_fd_sc_hd__o211a_1
X_11317_ hold4325/X _12365_/B _11316_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11317_/X
+ sky130_fd_sc_hd__o211a_1
X_15085_ _15193_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12297_ hold4656/X _13716_/A _12296_/X vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_201_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14036_ _15543_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_226_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11248_ hold3924/X _11726_/B _11247_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11248_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11179_ _11194_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _16883_/D sky130_fd_sc_hd__nor2_1
XTAP_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _16126_/CLK _15987_/D vssd1 vssd1 vccd1 vccd1 hold854/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _17726_/CLK _17726_/D vssd1 vssd1 vccd1 vccd1 _17726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14938_ _15207_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_380_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17742_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17657_ _17689_/CLK _17657_/D vssd1 vssd1 vccd1 vccd1 _17657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14869_ hold1710/X _14880_/B _14868_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16608_ _18228_/CLK _16608_/D vssd1 vssd1 vccd1 vccd1 _16608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08390_ _14894_/A hold1536/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_175_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _17642_/CLK _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16539_ _18223_/CLK _16539_/D vssd1 vssd1 vccd1 vccd1 _16539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _09053_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _16122_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18209_ _18209_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5804 output75/X vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5815 hold5951/X vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5826 _17525_/Q vssd1 vssd1 vccd1 vccd1 hold5826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 hold311/X vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 hold249/X vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5837 hold5974/X vssd1 vssd1 vccd1 vccd1 hold5837/X sky130_fd_sc_hd__clkbuf_2
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5848 hold5848/A vssd1 vssd1 vccd1 vccd1 hold5848/X sky130_fd_sc_hd__buf_2
Xhold5859 hold6018/X vssd1 vssd1 vccd1 vccd1 hold5859/X sky130_fd_sc_hd__clkbuf_4
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__clkbuf_16
Xhold145 hold5/X vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__buf_4
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09913_ hold4063/X _10007_/B _09912_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold178 la_data_in[18] vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _09366_/Y vssd1 vssd1 vccd1 vccd1 _09386_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout614 _09356_/Y vssd1 vssd1 vccd1 vccd1 _09357_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout625 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15481_/A1 sky130_fd_sc_hd__buf_4
Xfanout636 hold5900/X vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09844_ hold5054/X _10034_/B _09843_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09844_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout647 _13714_/C1 vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__buf_4
XFILLER_0_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout658 _12987_/A vssd1 vssd1 vccd1 vccd1 _12990_/A sky130_fd_sc_hd__buf_4
Xfanout669 fanout692/X vssd1 vssd1 vccd1 vccd1 _13801_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_241_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ hold4709/X _10577_/B _09774_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09775_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08726_ _09053_/A hold713/X vssd1 vssd1 vccd1 vccd1 _15984_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ hold292/X hold872/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ hold140/X hold335/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold336/A sky130_fd_sc_hd__mux2_1
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ hold1519/X hold3916/X _10997_/S vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ hold2882/X _09216_/B _09208_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09209_/X
+ sky130_fd_sc_hd__o211a_1
X_10481_ hold1718/X _16651_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ hold5296/X _12314_/B _12219_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _12220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_42_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_42_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_12151_ hold4417/X _12365_/B _12150_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ hold1634/X _16858_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__mux2_1
X_12082_ hold3478/X _12274_/A2 _12081_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12082_/X
+ sky130_fd_sc_hd__o211a_1
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__buf_6
XFILLER_0_120_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15910_ _16077_/CLK _15910_/D vssd1 vssd1 vccd1 vccd1 _15910_/Q sky130_fd_sc_hd__dfxtp_1
X_11033_ hold2701/X hold5044/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ _18032_/CLK _16890_/D vssd1 vssd1 vccd1 vccd1 _16890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _17732_/CLK _15841_/D vssd1 vssd1 vccd1 vccd1 _15841_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _08436_/X vssd1 vssd1 vccd1 vccd1 _15848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_138_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2091 _09135_/X vssd1 vssd1 vccd1 vccd1 _16180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _17721_/CLK _15772_/D vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfxtp_1
X_12984_ _12987_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _17504_/D sky130_fd_sc_hd__and2_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 _14901_/X vssd1 vssd1 vccd1 vccd1 _18236_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17517_/CLK _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14723_ hold2365/X _14714_/B _14722_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ hold5254/X _12314_/B _11934_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _15209_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14654_/X sky130_fd_sc_hd__or2_1
X_17442_ _17446_/CLK _17442_/D vssd1 vssd1 vccd1 vccd1 _17442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ hold4543/X _12344_/B _11865_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11866_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13713_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ hold2709/X hold5379/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14585_ hold2703/X _14612_/B _14584_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14585_/X
+ sky130_fd_sc_hd__o211a_1
X_17373_ _17376_/CLK _17373_/D vssd1 vssd1 vccd1 vccd1 _17373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _12367_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _17089_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16324_ _18375_/CLK _16324_/D vssd1 vssd1 vccd1 vccd1 _16324_/Q sky130_fd_sc_hd__dfxtp_1
X_13536_ _13767_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ _17941_/Q hold5463/X _11159_/C vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ _17378_/CLK _16255_/D vssd1 vssd1 vccd1 vccd1 _16255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13467_ _13788_/A _13467_/B vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ hold1658/X hold4666/X _11159_/C vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15206_ hold1092/X _15221_/B _15205_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15206_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12418_ _12418_/A _12418_/B vssd1 vssd1 vccd1 vccd1 _17302_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16186_ _17506_/CLK _16186_/D vssd1 vssd1 vccd1 vccd1 _16186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13398_ _13782_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__or2_1
X_15137_ _15191_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__or2_1
X_12349_ _13873_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _17273_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3709 _09589_/X vssd1 vssd1 vccd1 vccd1 _16353_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _15068_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _15068_/X sky130_fd_sc_hd__and2_1
XFILLER_0_227_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14019_ hold3071/X _14040_/B _14018_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _14019_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07890_ _14794_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07890_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ hold1581/X _13222_/A _10190_/S vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08511_ _15515_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17709_ _17741_/CLK _17709_/D vssd1 vssd1 vccd1 vccd1 _17709_/Q sky130_fd_sc_hd__dfxtp_1
X_09491_ _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13056_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_188_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ hold2420/X _08433_/B _08441_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _08442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ _08373_/A hold470/X vssd1 vssd1 vccd1 vccd1 _15818_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5601 _17011_/Q vssd1 vssd1 vccd1 vccd1 hold5601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5612 _10912_/X vssd1 vssd1 vccd1 vccd1 _16794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5623 _16951_/Q vssd1 vssd1 vccd1 vccd1 hold5623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5634 _10741_/X vssd1 vssd1 vccd1 vccd1 _16737_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4900 _10240_/X vssd1 vssd1 vccd1 vccd1 _16570_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5645 _16949_/Q vssd1 vssd1 vccd1 vccd1 hold5645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4911 _16716_/Q vssd1 vssd1 vccd1 vccd1 hold4911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5656 _10059_/Y vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4922 _10153_/X vssd1 vssd1 vccd1 vccd1 _16541_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5667 _17571_/Q vssd1 vssd1 vccd1 vccd1 hold5667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4933 _10513_/X vssd1 vssd1 vccd1 vccd1 _16661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5678 _09772_/X vssd1 vssd1 vccd1 vccd1 _16414_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4944 _16591_/Q vssd1 vssd1 vccd1 vccd1 hold4944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5689 _17599_/Q vssd1 vssd1 vccd1 vccd1 hold5689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4955 _10417_/X vssd1 vssd1 vccd1 vccd1 _16629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4966 _16997_/Q vssd1 vssd1 vccd1 vccd1 hold4966/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout400 _14393_/Y vssd1 vssd1 vccd1 vccd1 _14446_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4977 _11818_/X vssd1 vssd1 vccd1 vccd1 _17096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout411 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14202_/B sky130_fd_sc_hd__buf_6
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4988 _17692_/Q vssd1 vssd1 vccd1 vccd1 hold4988/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout422 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13995_/A2 sky130_fd_sc_hd__buf_8
Xhold4999 _11790_/Y vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout433 _13622_/S vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout444 _10025_/C vssd1 vssd1 vccd1 vccd1 _13622_/S sky130_fd_sc_hd__buf_4
Xfanout455 _11150_/C vssd1 vssd1 vccd1 vccd1 _11168_/C sky130_fd_sc_hd__clkbuf_4
Xfanout466 _10025_/C vssd1 vssd1 vccd1 vccd1 _13874_/C sky130_fd_sc_hd__clkbuf_8
X_09827_ _18344_/Q hold4036/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__mux2_1
Xfanout477 _11480_/S vssd1 vssd1 vccd1 vccd1 _12365_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_232_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout488 _10004_/C vssd1 vssd1 vccd1 vccd1 _10034_/C sky130_fd_sc_hd__buf_6
Xfanout499 _10400_/S vssd1 vssd1 vccd1 vccd1 _11096_/S sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_231_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16631_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_216_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ hold1194/X hold4843/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ hold607/X hold899/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold900/A sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ hold2146/X _16387_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__mux2_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _17064_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__and3_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ hold2132/X _17041_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ hold4636/X _10488_/A _10601_/X vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ _14370_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _17982_/D sky130_fd_sc_hd__and2_1
X_11582_ hold1668/X hold5501/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ hold4133/X _13814_/B _13320_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10533_ _10533_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16040_ _18410_/CLK _16040_/D vssd1 vssd1 vccd1 vccd1 hold672/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ hold3720/X _13251_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__mux2_2
X_10464_ _10560_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ hold2816/X _17225_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__mux2_1
X_13183_ _13199_/A1 _13181_/X _13182_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10395_ _10533_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12134_ hold1691/X hold4217/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17991_ _18059_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_319_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ hold2828/X hold5431/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__mux2_1
X_16942_ _17852_/CLK _16942_/D vssd1 vssd1 vccd1 vccd1 _16942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ _11124_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__or2_1
XFILLER_0_217_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16873_ _18042_/CLK _16873_/D vssd1 vssd1 vccd1 vccd1 _16873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15824_ _17639_/CLK _15824_/D vssd1 vssd1 vccd1 vccd1 _15824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ hold3065/X _17500_/Q _12967_/S vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__mux2_1
X_15755_ _17740_/CLK _15755_/D vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14706_ _15099_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__or2_1
X_11918_ hold1314/X hold4079/X _12302_/C vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__mux2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15686_ _17113_/CLK _15686_/D vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfxtp_1
X_12898_ hold2035/X hold3167/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux2_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17425_ _17425_/CLK _17425_/D vssd1 vssd1 vccd1 vccd1 _17425_/Q sky130_fd_sc_hd__dfxtp_1
X_14637_ hold2652/X _14664_/B _14636_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14637_/X
+ sky130_fd_sc_hd__o211a_1
X_11849_ hold2965/X hold4695/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11850_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ hold690/X _14573_/B hold2109/X vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__a21o_1
X_17356_ _17378_/CLK _17356_/D vssd1 vssd1 vccd1 vccd1 _17356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17815_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16307_ _16311_/CLK _16307_/D vssd1 vssd1 vccd1 vccd1 _16307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13519_ hold4166/X _13814_/B _13518_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13519_/X
+ sky130_fd_sc_hd__o211a_1
X_17287_ _17314_/CLK _17287_/D vssd1 vssd1 vccd1 vccd1 hold629/A sky130_fd_sc_hd__dfxtp_1
X_14499_ hold808/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16238_ _17420_/CLK _16238_/D vssd1 vssd1 vccd1 vccd1 _16238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4207 _17740_/Q vssd1 vssd1 vccd1 vccd1 hold4207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4218 _12040_/X vssd1 vssd1 vccd1 vccd1 _17170_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16169_ _17505_/CLK _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4229 _17234_/Q vssd1 vssd1 vccd1 vccd1 hold4229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3506 _17173_/Q vssd1 vssd1 vccd1 vccd1 hold3506/X sky130_fd_sc_hd__dlygate4sd3_1
X_08991_ hold140/X hold169/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__mux2_1
Xhold3517 _17647_/Q vssd1 vssd1 vccd1 vccd1 hold3517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3528 _12644_/X vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3539 _16351_/Q vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2805 _13993_/X vssd1 vssd1 vccd1 vccd1 _17801_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07942_ hold915/X _07986_/B vssd1 vssd1 vccd1 vccd1 _07942_/X sky130_fd_sc_hd__or2_1
Xhold2816 _15609_/Q vssd1 vssd1 vccd1 vccd1 hold2816/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2827 _14727_/X vssd1 vssd1 vccd1 vccd1 _18153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 _17901_/Q vssd1 vssd1 vccd1 vccd1 hold2838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2849 _09133_/X vssd1 vssd1 vccd1 vccd1 _16179_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07873_ _14330_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09612_ _09918_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09612_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09543_ _09963_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09474_ hold5910/X _09477_/C _09484_/B vssd1 vssd1 vccd1 vccd1 _09474_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08425_ _15213_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08356_ _15525_/A hold2999/X hold134/X vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08287_ hold915/X _08299_/B vssd1 vssd1 vccd1 vccd1 _08287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5420 _11932_/X vssd1 vssd1 vccd1 vccd1 _17134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5431 _17179_/Q vssd1 vssd1 vccd1 vccd1 hold5431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5442 _11668_/X vssd1 vssd1 vccd1 vccd1 _17046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5453 _16982_/Q vssd1 vssd1 vccd1 vccd1 hold5453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5464 _10654_/X vssd1 vssd1 vccd1 vccd1 _16708_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4730 _12354_/Y vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5475 _17053_/Q vssd1 vssd1 vccd1 vccd1 hold5475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4741 _16588_/Q vssd1 vssd1 vccd1 vccd1 hold4741/X sky130_fd_sc_hd__dlygate4sd3_1
X_10180_ hold4131/X _10598_/B _10179_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _10180_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5486 _10963_/X vssd1 vssd1 vccd1 vccd1 _16811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5497 _16980_/Q vssd1 vssd1 vccd1 vccd1 hold5497/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4752 _11733_/Y vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4763 _16407_/Q vssd1 vssd1 vccd1 vccd1 hold4763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4774 _10087_/X vssd1 vssd1 vccd1 vccd1 _16519_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_412_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4785 _16820_/Q vssd1 vssd1 vccd1 vccd1 hold4785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4796 _10561_/X vssd1 vssd1 vccd1 vccd1 _16677_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout230 _10622_/B vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__buf_4
XFILLER_0_234_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout241 _10037_/B vssd1 vssd1 vccd1 vccd1 _10477_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout252 _13698_/A vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout263 _11139_/A vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__buf_4
Xfanout274 _12231_/A vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__buf_4
Xfanout285 _11115_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__buf_4
XFILLER_0_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout296 _11061_/A vssd1 vssd1 vccd1 vccd1 _11136_/A sky130_fd_sc_hd__buf_4
XFILLER_0_195_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _13873_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _17743_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ hold3229/X _12820_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ hold2819/X _15547_/B _15539_/X _12657_/A vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__o211a_1
X_12752_ hold3414/X _12751_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__mux2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11703_ _12057_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__or2_1
X_15471_ _15489_/A _15471_/B _15471_/C _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_210_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ hold3756/X _12682_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17210_/CLK _17210_/D vssd1 vssd1 vccd1 vccd1 _17210_/Q sky130_fd_sc_hd__dfxtp_1
X_14422_ hold1863/X _14433_/B _14421_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _14422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11634_ _11637_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__or2_1
X_18190_ _18222_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14353_ _14910_/A hold2818/X hold333/X vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__mux2_1
X_17141_ _17153_/CLK _17141_/D vssd1 vssd1 vccd1 vccd1 _17141_/Q sky130_fd_sc_hd__dfxtp_1
X_11565_ _11667_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13297_/X _13303_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10516_ hold3980/X _10646_/B _10515_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17072_ _17886_/CLK _17072_/D vssd1 vssd1 vccd1 vccd1 _17072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14284_ hold808/A _14284_/B vssd1 vssd1 vccd1 vccd1 hold602/A sky130_fd_sc_hd__or2_1
XFILLER_0_165_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11496_ _12234_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ _17321_/CLK _16023_/D vssd1 vssd1 vccd1 vccd1 hold337/A sky130_fd_sc_hd__dfxtp_1
X_13235_ _13234_/X _16922_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__mux2_1
X_10447_ hold4986/X _10631_/B _10446_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _10447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _13166_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10378_ hold5182/X _10625_/B _10377_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_153_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16128_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12117_ _13797_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13097_ _13097_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__and2_1
X_17974_ _18038_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12048_ _12273_/A _12048_/B vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__or2_1
X_16925_ _17890_/CLK _16925_/D vssd1 vssd1 vccd1 vccd1 _16925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16856_ _18200_/CLK _16856_/D vssd1 vssd1 vccd1 vccd1 _16856_/Q sky130_fd_sc_hd__dfxtp_1
X_15807_ _17686_/CLK _15807_/D vssd1 vssd1 vccd1 vccd1 _15807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16787_ _17996_/CLK _16787_/D vssd1 vssd1 vccd1 vccd1 _16787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13999_ hold1624/X _13986_/B _13998_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _13999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _17741_/CLK _15738_/D vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _18460_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
X_15669_ _18428_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ hold2051/X _08209_/B _08209_/Y _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17408_ _18456_/CLK _17408_/D vssd1 vssd1 vccd1 vccd1 _17408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09190_ _15519_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18388_ _18394_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08141_ _08143_/A hold109/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__and2_1
X_17339_ _17339_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 _17339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08072_ _15531_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4004 hold5853/X vssd1 vssd1 vccd1 vccd1 hold5854/A sky130_fd_sc_hd__buf_4
XFILLER_0_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4015 _11629_/X vssd1 vssd1 vccd1 vccd1 _17033_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4026 _16452_/Q vssd1 vssd1 vccd1 vccd1 hold4026/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4037 _09733_/X vssd1 vssd1 vccd1 vccd1 _16401_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4048 _16975_/Q vssd1 vssd1 vccd1 vccd1 hold4048/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3303 _17466_/Q vssd1 vssd1 vccd1 vccd1 hold3303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4059 _16424_/Q vssd1 vssd1 vccd1 vccd1 hold4059/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3314 _17463_/Q vssd1 vssd1 vccd1 vccd1 hold3314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3325 _17465_/Q vssd1 vssd1 vccd1 vccd1 hold3325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3336 _17388_/Q vssd1 vssd1 vccd1 vccd1 hold3336/X sky130_fd_sc_hd__dlygate4sd3_1
X_08974_ _12438_/A hold481/X vssd1 vssd1 vccd1 vccd1 _16104_/D sky130_fd_sc_hd__and2_1
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2602 _08057_/X vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3347 _17440_/Q vssd1 vssd1 vccd1 vccd1 hold3347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3358 _09709_/X vssd1 vssd1 vccd1 vccd1 _16393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _08089_/X vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3369 _09793_/X vssd1 vssd1 vccd1 vccd1 _16421_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2624 _17902_/Q vssd1 vssd1 vccd1 vccd1 hold2624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _14472_/X vssd1 vssd1 vccd1 vccd1 _18031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 _18022_/Q vssd1 vssd1 vccd1 vccd1 hold1901/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ hold2302/X _07924_/B _07924_/Y _08163_/A vssd1 vssd1 vccd1 vccd1 _07925_/X
+ sky130_fd_sc_hd__o211a_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_1
Xhold2646 _07947_/X vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1912 _18133_/Q vssd1 vssd1 vccd1 vccd1 hold1912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 _08032_/X vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _18234_/Q vssd1 vssd1 vccd1 vccd1 hold1923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _07915_/X vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _14845_/X vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 _18247_/Q vssd1 vssd1 vccd1 vccd1 hold2679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1945 _18164_/Q vssd1 vssd1 vccd1 vccd1 hold1945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1956 _18086_/Q vssd1 vssd1 vccd1 vccd1 hold1956/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ hold2780/X _07869_/B _07855_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07856_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1967 _15005_/X vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1978 _14861_/X vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _14325_/X vssd1 vssd1 vccd1 vccd1 _17960_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _12310_/A vssd1 vssd1 vccd1 vccd1 _07787_/Y sky130_fd_sc_hd__inv_4
XFILLER_0_17_1310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ hold3808/X _10004_/B _09525_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09463_/D _09484_/B _09457_/C vssd1 vssd1 vccd1 vccd1 _16312_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ hold2174/X _08440_/A2 _08407_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _08408_/X
+ sky130_fd_sc_hd__o211a_1
X_09388_ hold5844/A _09342_/B _09342_/Y _09387_/X _12404_/A vssd1 vssd1 vccd1 vccd1
+ _09388_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08339_ hold203/A hold331/A vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__or2_1
XFILLER_0_145_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ hold5449/X _11732_/B _11349_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10301_ hold1642/X _16591_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ hold5645/X _11768_/B _11280_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _11281_/X
+ sky130_fd_sc_hd__o211a_1
X_13020_ _09489_/B hold954/X vssd1 vssd1 vccd1 vccd1 hold955/A sky130_fd_sc_hd__nand2b_1
Xhold5250 _16974_/Q vssd1 vssd1 vccd1 vccd1 hold5250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5261 _10120_/X vssd1 vssd1 vccd1 vccd1 _16530_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10232_ hold2687/X hold3839/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__mux2_1
Xhold5272 _17232_/Q vssd1 vssd1 vccd1 vccd1 hold5272/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5283 _13480_/X vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5294 _17041_/Q vssd1 vssd1 vccd1 vccd1 hold5294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4560 _13549_/X vssd1 vssd1 vccd1 vccd1 _17636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4571 _16004_/Q vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10163_ hold2830/X hold3575/X _10997_/S vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__mux2_1
Xhold4582 _15443_/X vssd1 vssd1 vccd1 vccd1 _15444_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4593 hold5875/X vssd1 vssd1 vccd1 vccd1 hold5876/A sky130_fd_sc_hd__buf_4
XFILLER_0_238_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3870 _17066_/Q vssd1 vssd1 vccd1 vccd1 hold3870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3881 _09547_/X vssd1 vssd1 vccd1 vccd1 _16339_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14971_ hold1678/X hold514/X _14970_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14971_/X
+ sky130_fd_sc_hd__o211a_1
X_10094_ hold2120/X hold4606/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__mux2_1
Xhold3892 _16577_/Q vssd1 vssd1 vccd1 vccd1 hold3892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16710_ _18039_/CLK _16710_/D vssd1 vssd1 vccd1 vccd1 _16710_/Q sky130_fd_sc_hd__dfxtp_1
X_13922_ _15211_/A _17767_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 _13922_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17690_ _17722_/CLK _17690_/D vssd1 vssd1 vccd1 vccd1 _17690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _18229_/CLK _16641_/D vssd1 vssd1 vccd1 vccd1 _16641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13853_ _17738_/Q _13886_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__and3_1
XFILLER_0_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ _12804_/A _12804_/B vssd1 vssd1 vccd1 vccd1 _17444_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16572_ _18180_/CLK _16572_/D vssd1 vssd1 vccd1 vccd1 _16572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ hold5166/X _11198_/B _10995_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10996_/X
+ sky130_fd_sc_hd__o211a_1
X_13784_ hold2359/X hold4374/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18311_ _18331_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__dfxtp_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _15523_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12738_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _17421_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_1307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18396_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15454_/A _15454_/B vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__and2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12759_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _17398_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ hold3784/X _11617_/A2 _11616_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _17029_/D
+ sky130_fd_sc_hd__o211a_1
X_14405_ _15193_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__or2_1
X_18173_ _18201_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_6_1_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_15385_ _15385_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__or2_1
X_12597_ _12600_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _17375_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ _17188_/CLK _17124_/D vssd1 vssd1 vccd1 vccd1 _17124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ hold5270/X _11738_/B _11547_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11548_/X
+ sky130_fd_sc_hd__o211a_1
X_14336_ _14443_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_334_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold519 hold519/A vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ hold2351/X _14266_/B _14266_/Y _15194_/C1 vssd1 vssd1 vccd1 vccd1 _14267_/X
+ sky130_fd_sc_hd__o211a_1
X_17055_ _17891_/CLK _17055_/D vssd1 vssd1 vccd1 vccd1 _17055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ hold5647/X _11789_/B _11478_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _16983_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16006_ _18411_/CLK _16006_/D vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _17578_/Q _17112_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14198_ _14878_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_221_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13148_/X hold3553/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17957_ _18053_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _17812_/Q vssd1 vssd1 vccd1 vccd1 hold1208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _14558_/X vssd1 vssd1 vccd1 vccd1 hold1219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ _17822_/CLK _16908_/D vssd1 vssd1 vccd1 vccd1 _16908_/Q sky130_fd_sc_hd__dfxtp_1
X_08690_ _12416_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _15966_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17888_ _17888_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16839_ _18040_/CLK _16839_/D vssd1 vssd1 vccd1 vccd1 _16839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18071_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_221_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _15099_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ _12768_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _16232_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ hold2832/X _09177_/A2 _09172_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08124_ _15529_/A hold2572/X hold240/X vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08055_ hold2616/X _08097_/A2 _08054_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _08055_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3100 _16262_/Q vssd1 vssd1 vccd1 vccd1 hold3100/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3111 _14317_/X vssd1 vssd1 vccd1 vccd1 _17956_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3122 _18165_/Q vssd1 vssd1 vccd1 vccd1 hold3122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3133 _14466_/X vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3144 _14755_/X vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2410 _14079_/X vssd1 vssd1 vccd1 vccd1 _17842_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3155 _17356_/Q vssd1 vssd1 vccd1 vccd1 hold3155/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3166 _14253_/X vssd1 vssd1 vccd1 vccd1 _17925_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2421 _08442_/X vssd1 vssd1 vccd1 vccd1 _15851_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3177 _17441_/Q vssd1 vssd1 vccd1 vccd1 hold3177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 _17935_/Q vssd1 vssd1 vccd1 vccd1 hold2432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2443 _18213_/Q vssd1 vssd1 vccd1 vccd1 hold2443/X sky130_fd_sc_hd__dlygate4sd3_1
X_08957_ hold361/X hold783/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold784/A sky130_fd_sc_hd__mux2_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3188 _12818_/X vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2454 _14231_/X vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1720 _17937_/Q vssd1 vssd1 vccd1 vccd1 hold1720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3199 _17423_/Q vssd1 vssd1 vccd1 vccd1 hold3199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2465 _18168_/Q vssd1 vssd1 vccd1 vccd1 hold2465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1731 _18131_/Q vssd1 vssd1 vccd1 vccd1 hold1731/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2476 _08510_/X vssd1 vssd1 vccd1 vccd1 _15882_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07908_ _14758_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08888_ hold163/X hold314/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold315/A sky130_fd_sc_hd__mux2_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1742 _15764_/Q vssd1 vssd1 vccd1 vccd1 hold1742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2487 _08040_/X vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2498 _18116_/Q vssd1 vssd1 vccd1 vccd1 hold2498/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1753 _17943_/Q vssd1 vssd1 vccd1 vccd1 hold1753/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1764 _14139_/X vssd1 vssd1 vccd1 vccd1 _17871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 _16162_/Q vssd1 vssd1 vccd1 vccd1 hold1775/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _14403_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1786 _08046_/X vssd1 vssd1 vccd1 vccd1 _15664_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1797 _18092_/Q vssd1 vssd1 vccd1 vccd1 hold1797/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ hold1476/X _16774_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_196_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _18238_/Q _13086_/A _10019_/C vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__mux2_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ hold2921/X _16751_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _10782_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_195_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ hold1404/X _17351_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ hold215/X _12509_/A2 _12507_/A3 _12450_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold96/A sky130_fd_sc_hd__o311a_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11402_ hold1624/X _16958_/Q _11594_/S vssd1 vssd1 vccd1 vccd1 _11403_/B sky130_fd_sc_hd__mux2_1
X_15170_ hold2284/X _15165_/B _15169_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _15170_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12382_ _12531_/A hold705/X vssd1 vssd1 vccd1 vccd1 _17284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_90 hold746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14121_ hold1650/X _14142_/B _14120_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ hold2888/X hold5014/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _15233_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ hold1348/X hold3567/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11265_/B sky130_fd_sc_hd__mux2_1
X_13003_ _14897_/A hold533/X vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__nor2_2
Xhold5080 _17596_/Q vssd1 vssd1 vccd1 vccd1 hold5080/X sky130_fd_sc_hd__dlygate4sd3_1
X_10215_ _10563_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__or2_1
Xhold5091 _09868_/X vssd1 vssd1 vccd1 vccd1 _16446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195_ _16889_/Q _11762_/B _11762_/C vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4390 _13396_/X vssd1 vssd1 vccd1 vccd1 _17585_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17811_ _18425_/CLK _17811_/D vssd1 vssd1 vccd1 vccd1 _17811_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10146_ _10476_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2_1
XTAP_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17742_ _17742_/CLK _17742_/D vssd1 vssd1 vccd1 vccd1 _17742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14954_ hold972/X _14958_/B vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__or2_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ _10563_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10077_/X sky130_fd_sc_hd__or2_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ _13905_/A _13905_/B vssd1 vssd1 vccd1 vccd1 _17758_/D sky130_fd_sc_hd__and2_1
X_17673_ _17737_/CLK _17673_/D vssd1 vssd1 vccd1 vccd1 _17673_/Q sky130_fd_sc_hd__dfxtp_1
X_14885_ hold1001/X _14882_/B _14884_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14885_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ _18186_/CLK _16624_/D vssd1 vssd1 vccd1 vccd1 _16624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ hold3988/X _13761_/A _13835_/X vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16555_ _18175_/CLK _16555_/D vssd1 vssd1 vccd1 vccd1 _16555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10979_ hold1406/X hold3926/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__mux2_1
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15506_ _15506_/A _15506_/B vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__and2_1
X_12718_ _16237_/Q hold3372/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _18397_/CLK _16486_/D vssd1 vssd1 vccd1 vccd1 _16486_/Q sky130_fd_sc_hd__dfxtp_1
X_13698_ _13698_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__or2_1
X_18225_ _18225_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
X_15437_ hold783/X _09392_/B _09392_/C hold652/X vssd1 vssd1 vccd1 vccd1 _15437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ hold2782/X _17394_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18156_ _18220_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15368_ hold286/X _15484_/A2 _09392_/D hold508/X vssd1 vssd1 vccd1 vccd1 _15368_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ _17899_/CLK _17107_/D vssd1 vssd1 vccd1 vccd1 _17107_/Q sky130_fd_sc_hd__dfxtp_1
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14319_ hold2753/X _14326_/B _14318_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14319_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18087_ _18175_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15299_ hold789/X _15485_/A2 _15488_/A2 hold862/X _15298_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold327 hold686/X vssd1 vssd1 vccd1 vccd1 hold687/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17038_ _17884_/CLK _17038_/D vssd1 vssd1 vccd1 vccd1 _17038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09860_ hold3134/X _16444_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__mux2_1
Xfanout807 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _15222_/C1 sky130_fd_sc_hd__buf_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout818 _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15162_/C1 sky130_fd_sc_hd__buf_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout829 _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14542_/C1 sky130_fd_sc_hd__buf_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _09061_/A hold252/X vssd1 vssd1 vccd1 vccd1 _16024_/D sky130_fd_sc_hd__and2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ hold2963/X _16421_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _18303_/Q vssd1 vssd1 vccd1 vccd1 hold1005/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1016 _15535_/A vssd1 vssd1 vccd1 vccd1 hold1016/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _15364_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__and2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _09071_/X vssd1 vssd1 vccd1 vccd1 _16150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 _17913_/Q vssd1 vssd1 vccd1 vccd1 hold1038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _15152_/X vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08673_ hold88/X hold127/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_206_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_256_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18124_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09225_ hold2808/X _09216_/B _09224_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _09225_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09156_ _15539_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08107_ _15498_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _15692_/D sky130_fd_sc_hd__and2_1
Xclkbuf_6_32_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_32_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09087_ hold968/X _09119_/A2 _09086_/X _12987_/A vssd1 vssd1 vccd1 vccd1 hold969/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08038_ hold1258/X _08033_/B _08037_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _08038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold850 hold850/A vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold861 hold861/A vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold872 hold872/A vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 hold894/A vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _11158_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _16490_/D sky130_fd_sc_hd__nor2_1
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _16487_/Q _10013_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__and3_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 _17863_/Q vssd1 vssd1 vccd1 vccd1 hold2240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 _15192_/X vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2262 _18014_/Q vssd1 vssd1 vccd1 vccd1 hold2262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2273 _18314_/Q vssd1 vssd1 vccd1 vccd1 hold2273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2284 _18366_/Q vssd1 vssd1 vccd1 vccd1 hold2284/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2295 _15844_/Q vssd1 vssd1 vccd1 vccd1 hold2295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 _14045_/X vssd1 vssd1 vccd1 vccd1 _17826_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1561 _17831_/Q vssd1 vssd1 vccd1 vccd1 hold1561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1572 _15150_/X vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ hold2424/X _17141_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__mux2_1
Xhold1583 _16256_/Q vssd1 vssd1 vccd1 vccd1 hold1583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1594 _14235_/X vssd1 vssd1 vccd1 vccd1 _17916_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ _10998_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14670_ _15225_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__or2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _15710_/Q hold3623/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ _11121_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10833_/X sky130_fd_sc_hd__or2_1
X_13621_ hold4988/X _13811_/B _13620_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _18321_/CLK _16340_/D vssd1 vssd1 vccd1 vccd1 _16340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _11052_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13552_ hold4358/X _13856_/B _13551_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ hold11/X _12445_/A _12445_/B _12502_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold12/A sky130_fd_sc_hd__o311a_1
XFILLER_0_164_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16271_ _17376_/CLK _16271_/D vssd1 vssd1 vccd1 vccd1 _16271_/Q sky130_fd_sc_hd__dfxtp_1
X_13483_ hold5737/X _13817_/B _13482_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _13483_/X
+ sky130_fd_sc_hd__o211a_1
X_10695_ _11115_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _18010_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ _13037_/A hold323/X vssd1 vssd1 vccd1 vccd1 _17310_/D sky130_fd_sc_hd__and2_1
X_15222_ hold1493/X _15221_/B _15221_/Y _15222_/C1 vssd1 vssd1 vccd1 vccd1 _15222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15153_ _15207_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15153_/X sky130_fd_sc_hd__or2_1
X_12365_ _12365_/A _12365_/B _12365_/C vssd1 vssd1 vccd1 vccd1 _12365_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11316_ _12246_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__or2_1
X_14104_ _14443_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ hold2208/X _15111_/B _15083_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15084_/X
+ sky130_fd_sc_hd__o211a_1
X_12296_ _17256_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ hold2426/X _14040_/B _14034_/Y _13927_/A vssd1 vssd1 vccd1 vccd1 _14035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _11631_/A _11247_/B vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11178_ hold4664/X _11082_/A _11177_/X vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_219_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10129_ hold4958/X _10631_/B _10128_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ _16131_/CLK _15986_/D vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__dfxtp_1
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _17725_/CLK _17725_/D vssd1 vssd1 vccd1 vccd1 _17725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14937_ hold1273/X _14952_/B _14936_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14937_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17656_ _17726_/CLK _17656_/D vssd1 vssd1 vccd1 vccd1 _17656_/Q sky130_fd_sc_hd__dfxtp_1
X_14868_ _15207_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16607_ _18131_/CLK _16607_/D vssd1 vssd1 vccd1 vccd1 _16607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13819_ _13825_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _17726_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_159_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17587_ _17683_/CLK _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
X_14799_ hold2216/X _14826_/B _14798_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14799_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16538_ _18222_/CLK _16538_/D vssd1 vssd1 vccd1 vccd1 _16538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _18316_/CLK _16469_/D vssd1 vssd1 vccd1 vccd1 _16469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ hold17/X hold224/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ _18208_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5805 hold5942/X vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__buf_1
X_18139_ _18205_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5816 output72/X vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_223_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5827 _17519_/Q vssd1 vssd1 vccd1 vccd1 hold5827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold251/X vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__clkbuf_4
Xhold5838 hold5838/A vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_12
Xhold5849 hold6010/X vssd1 vssd1 vccd1 vccd1 hold5849/X sky130_fd_sc_hd__buf_2
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__buf_12
XFILLER_0_223_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _09936_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__or2_1
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 input46/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout604 _09364_/Y vssd1 vssd1 vccd1 vccd1 _09392_/D sky130_fd_sc_hd__buf_6
XFILLER_0_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout615 _09356_/Y vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__clkbuf_4
Xfanout626 hold202/X vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__clkbuf_2
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__or2_1
Xfanout637 _12696_/A vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__clkbuf_4
Xfanout648 fanout693/X vssd1 vssd1 vccd1 vccd1 _13714_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout659 fanout693/X vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__buf_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09774_ _10482_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__or2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ hold498/X hold712/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold713/A sky130_fd_sc_hd__mux2_1
XFILLER_0_241_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _12408_/A hold287/X vssd1 vssd1 vccd1 vccd1 _15950_/D sky130_fd_sc_hd__and2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_437_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17726_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08587_ _15414_/A hold159/X vssd1 vssd1 vccd1 vccd1 _15917_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _15537_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ hold4745/X _11192_/B _10479_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09139_ hold2096/X _09177_/A2 _09138_/X _12912_/A vssd1 vssd1 vccd1 vccd1 _09139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12150_ _12246_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11101_ hold4893/X _11180_/B _11100_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11101_/X
+ sky130_fd_sc_hd__o211a_1
X_12081_ _13782_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__or2_1
Xhold680 hold680/A vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold691 hold691/A vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__buf_4
XFILLER_0_229_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ hold5643/X _11207_/B _11031_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _11032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15840_ _17244_/CLK _15840_/D vssd1 vssd1 vccd1 vccd1 _15840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _15787_/Q vssd1 vssd1 vccd1 vccd1 hold2070/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2081 _18435_/Q vssd1 vssd1 vccd1 vccd1 hold2081/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 _17962_/Q vssd1 vssd1 vccd1 vccd1 hold2092/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _17426_/CLK _15771_/D vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ hold3138/X _12982_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_232_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17510_/CLK _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1380 _08340_/X vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ _15169_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__or2_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1391 _17852_/Q vssd1 vssd1 vccd1 vccd1 hold1391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _12219_/A _11934_/B vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__or2_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17446_/CLK _17441_/D vssd1 vssd1 vccd1 vccd1 _17441_/Q sky130_fd_sc_hd__dfxtp_1
X_14653_ hold3055/X _14664_/B _14652_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14653_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _12057_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17297_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13604_ hold2836/X hold3938/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__mux2_1
X_17372_ _17372_/CLK _17372_/D vssd1 vssd1 vccd1 vccd1 _17372_/Q sky130_fd_sc_hd__dfxtp_1
X_10816_ hold4419/X _11207_/B _10815_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10816_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14584_ _15193_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14584_/X sky130_fd_sc_hd__or2_1
X_11796_ hold3670/X _12246_/A _11795_/X vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16323_ _16323_/CLK _16323_/D vssd1 vssd1 vccd1 vccd1 _16323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ hold2537/X _17632_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ hold5573/X _11789_/B _10746_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _10747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ _17378_/CLK _16254_/D vssd1 vssd1 vccd1 vccd1 _16254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10678_ hold5300/X _11159_/B _10677_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _10678_/X
+ sky130_fd_sc_hd__o211a_1
X_13466_ hold1929/X _17609_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13467_/B sky130_fd_sc_hd__mux2_1
X_15205_ _15205_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__or2_1
X_12417_ hold568/X hold792/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12418_/B sky130_fd_sc_hd__mux2_1
X_16185_ _17506_/CLK hold976/X vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ hold1538/X hold3740/X _13877_/C vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ hold3139/X _15167_/B _15135_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _15136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ hold3596/X _13773_/A _12347_/X vssd1 vssd1 vccd1 vccd1 _12348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15067_ _15121_/A _18317_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__mux2_1
X_12279_ _13461_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14018_ _15525_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15969_ _16077_/CLK _15969_/D vssd1 vssd1 vccd1 vccd1 hold374/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ hold2475/X _08503_/Y _08509_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17708_ _17740_/CLK _17708_/D vssd1 vssd1 vccd1 vccd1 _17708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ _13029_/A _13043_/C hold990/X vssd1 vssd1 vccd1 vccd1 _13055_/C sky130_fd_sc_hd__and3_4
XFILLER_0_210_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08441_ _14782_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _17639_/CLK _17639_/D vssd1 vssd1 vccd1 vccd1 _17639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ hold469/X _15818_/Q hold134/X vssd1 vssd1 vccd1 vccd1 hold470/A sky130_fd_sc_hd__mux2_1
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5602 _11467_/X vssd1 vssd1 vccd1 vccd1 _16979_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5613 _17087_/Q vssd1 vssd1 vccd1 vccd1 hold5613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5624 _11287_/X vssd1 vssd1 vccd1 vccd1 _16919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5635 _16859_/Q vssd1 vssd1 vccd1 vccd1 hold5635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4901 _16552_/Q vssd1 vssd1 vccd1 vccd1 hold4901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5646 _11281_/X vssd1 vssd1 vccd1 vccd1 _16917_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4912 _11157_/Y vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5657 _17570_/Q vssd1 vssd1 vccd1 vccd1 hold5657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4923 _16707_/Q vssd1 vssd1 vccd1 vccd1 hold4923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5668 _13833_/Y vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4934 _17630_/Q vssd1 vssd1 vccd1 vccd1 hold4934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5679 _16414_/Q vssd1 vssd1 vccd1 vccd1 hold5679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4945 _10207_/X vssd1 vssd1 vccd1 vccd1 _16559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4956 _17256_/Q vssd1 vssd1 vccd1 vccd1 hold4956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4967 _11425_/X vssd1 vssd1 vccd1 vccd1 _16965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4978 _16643_/Q vssd1 vssd1 vccd1 vccd1 hold4978/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout401 hold332/X vssd1 vssd1 vccd1 vccd1 hold333/A sky130_fd_sc_hd__buf_6
Xfanout412 _14140_/B vssd1 vssd1 vccd1 vccd1 _14160_/B sky130_fd_sc_hd__buf_8
XFILLER_0_217_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4989 _13621_/X vssd1 vssd1 vccd1 vccd1 _17660_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout423 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__clkbuf_8
Xfanout434 _12302_/C vssd1 vssd1 vccd1 vccd1 _13811_/C sky130_fd_sc_hd__clkbuf_8
Xfanout445 _11711_/S vssd1 vssd1 vccd1 vccd1 _12299_/C sky130_fd_sc_hd__clkbuf_8
Xfanout456 _10025_/C vssd1 vssd1 vccd1 vccd1 _11150_/C sky130_fd_sc_hd__buf_4
X_09826_ hold4473/X _09832_/A2 _09825_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _09826_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout467 _12368_/C vssd1 vssd1 vccd1 vccd1 _13556_/S sky130_fd_sc_hd__clkbuf_8
Xfanout478 _11480_/S vssd1 vssd1 vccd1 vccd1 _11792_/C sky130_fd_sc_hd__clkbuf_4
Xfanout489 _11057_/S vssd1 vssd1 vccd1 vccd1 _10004_/C sky130_fd_sc_hd__buf_6
X_09757_ hold3782/X _10007_/B _09756_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09757_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_240_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _12396_/A hold703/X vssd1 vssd1 vccd1 vccd1 _15975_/D sky130_fd_sc_hd__and2_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ hold5683/X _10070_/B _09687_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09688_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_271_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ hold353/X hold491/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_200_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ hold5174/X _12317_/B _11649_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11650_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10601_ _10601_/A _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__and3_1
X_11581_ hold4350/X _12338_/B _11580_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11581_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ hold1914/X hold4853/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__mux2_1
X_13320_ _13800_/A _13320_/B vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10463_ hold2002/X hold4028/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__mux2_1
X_13251_ _13250_/X _16924_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ hold4956/X _13811_/B _12201_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _12202_/X
+ sky130_fd_sc_hd__o211a_1
X_13182_ _13182_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__or2_1
X_10394_ hold1859/X _16622_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12133_ hold4305/X _13871_/B _12132_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _18229_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ hold4177/X _13868_/B _12063_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _12064_/X
+ sky130_fd_sc_hd__o211a_1
X_16941_ _17851_/CLK _16941_/D vssd1 vssd1 vccd1 vccd1 _16941_/Q sky130_fd_sc_hd__dfxtp_1
X_11015_ hold3031/X hold4425/X _11219_/C vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16872_ _18041_/CLK _16872_/D vssd1 vssd1 vccd1 vccd1 _16872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _17702_/CLK _15823_/D vssd1 vssd1 vccd1 vccd1 _15823_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_359_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17236_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _17641_/CLK _15754_/D vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _12969_/A _12966_/B vssd1 vssd1 vccd1 vccd1 _17498_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ hold2520/X _14720_/B _14704_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11917_ hold5248/X _12299_/B _11916_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _17113_/CLK _15685_/D vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12897_ _15502_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _17475_/D sky130_fd_sc_hd__and2_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _17426_/CLK _17424_/D vssd1 vssd1 vccd1 vccd1 _17424_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _15191_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14636_/X sky130_fd_sc_hd__or2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11848_ hold4261/X _13871_/B _11847_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _11848_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17355_ _17378_/CLK _17355_/D vssd1 vssd1 vccd1 vccd1 _17355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ _15191_/A _14557_/Y hold2007/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _14567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11779_ _13864_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _17083_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ _16311_/CLK _16306_/D vssd1 vssd1 vccd1 vccd1 _16306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _13713_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/X sky130_fd_sc_hd__or2_1
X_17286_ _17286_/CLK _17286_/D vssd1 vssd1 vccd1 vccd1 hold407/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14498_ hold1968/X _14487_/B _14497_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16237_ _17420_/CLK hold946/X vssd1 vssd1 vccd1 vccd1 _16237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13449_ _13698_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13449_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_75_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18010_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4208 _13765_/X vssd1 vssd1 vccd1 vccd1 _17708_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _17505_/CLK _16168_/D vssd1 vssd1 vccd1 vccd1 _16168_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4219 _16870_/Q vssd1 vssd1 vccd1 vccd1 hold4219/X sky130_fd_sc_hd__dlygate4sd3_1
X_15119_ _15227_/A hold734/X vssd1 vssd1 vccd1 vccd1 _15119_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3507 _11953_/X vssd1 vssd1 vccd1 vccd1 _17141_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16099_ _17322_/CLK _16099_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
X_08990_ _12436_/A hold197/X vssd1 vssd1 vccd1 vccd1 _16112_/D sky130_fd_sc_hd__and2_1
Xhold3518 _13486_/X vssd1 vssd1 vccd1 vccd1 _17615_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3529 _17608_/Q vssd1 vssd1 vccd1 vccd1 hold3529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07941_ hold1489/X _07991_/A2 _07940_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07941_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2806 _16188_/Q vssd1 vssd1 vccd1 vccd1 hold2806/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2817 _07931_/X vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 _15615_/Q vssd1 vssd1 vccd1 vccd1 hold2828/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2839 _14201_/X vssd1 vssd1 vccd1 vccd1 _17901_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ hold2363/X _07869_/B _07871_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07872_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09611_ _18272_/Q hold3361/X _10019_/C vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_223_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ hold1672/X _13174_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _09477_/C _09484_/B _09473_/C vssd1 vssd1 vccd1 vccd1 _16318_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08424_ hold5991/X _08433_/B hold1357/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08424_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08355_ _12747_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _15809_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ hold1340/X _08336_/A2 _08285_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5410 _10882_/X vssd1 vssd1 vccd1 vccd1 _16784_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5421 _17276_/Q vssd1 vssd1 vccd1 vccd1 hold5421/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5432 _11971_/X vssd1 vssd1 vccd1 vccd1 _17147_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5443 _17148_/Q vssd1 vssd1 vccd1 vccd1 hold5443/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5454 _11380_/X vssd1 vssd1 vccd1 vccd1 _16950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4720 _12321_/Y vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5465 _17180_/Q vssd1 vssd1 vccd1 vccd1 hold5465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4731 _16384_/Q vssd1 vssd1 vccd1 vccd1 hold4731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5476 _11593_/X vssd1 vssd1 vccd1 vccd1 _17021_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4742 _10198_/X vssd1 vssd1 vccd1 vccd1 _16556_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5487 _16805_/Q vssd1 vssd1 vccd1 vccd1 hold5487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4753 _16788_/Q vssd1 vssd1 vccd1 vccd1 hold4753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5498 _11374_/X vssd1 vssd1 vccd1 vccd1 _16948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4764 _09655_/X vssd1 vssd1 vccd1 vccd1 _16375_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4775 _16549_/Q vssd1 vssd1 vccd1 vccd1 hold4775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4786 _10894_/X vssd1 vssd1 vccd1 vccd1 _16788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout220 fanout246/X vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__buf_8
Xhold4797 _16509_/Q vssd1 vssd1 vccd1 vccd1 hold4797/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout231 _10622_/B vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__buf_4
XFILLER_0_121_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout242 _10637_/B vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__buf_4
XFILLER_0_227_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout253 _13698_/A vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout264 _11652_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__buf_4
Xfanout275 _12231_/A vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__buf_4
XFILLER_0_226_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout286 _11115_/A vssd1 vssd1 vccd1 vccd1 _11667_/A sky130_fd_sc_hd__buf_4
X_09809_ hold885/X _16427_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__mux2_1
Xfanout297 _11061_/A vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_452_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ hold2027/X hold3184/X _12826_/S vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12751_ hold2178/X hold3403/X _12751_/S vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__mux2_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ hold1654/X _17058_/Q _12344_/C vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__mux2_1
X_15470_ hold708/X _09392_/C _15467_/X vssd1 vssd1 vccd1 vccd1 _15471_/D sky130_fd_sc_hd__a21o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12682_ hold2913/X _17405_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__mux2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14421_ _15535_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__or2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ hold1861/X _17035_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _17236_/CLK _17140_/D vssd1 vssd1 vccd1 vccd1 _17140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ _15496_/A hold487/X vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__and2_1
XFILLER_0_181_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ hold1446/X hold5513/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13303_ _13052_/X _13301_/X _13302_/X _13049_/Y vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_29_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ _10998_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17071_ _17834_/CLK _17071_/D vssd1 vssd1 vccd1 vccd1 _17071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14283_ hold1503/X _14272_/B _14282_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _14283_/X
+ sky130_fd_sc_hd__o211a_1
X_11495_ hold2236/X _16989_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16022_ _17347_/CLK _16022_/D vssd1 vssd1 vccd1 vccd1 _16022_/Q sky130_fd_sc_hd__dfxtp_1
X_10446_ _10542_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13234_ _17580_/Q _17114_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13165_ _13164_/X hold4725/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__mux2_1
X_10377_ _10560_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ hold2269/X _17196_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__mux2_1
X_13096_ _13089_/X _13095_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17530_/D sky130_fd_sc_hd__o21a_1
X_17973_ _18071_/CLK hold488/X vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12047_ hold2486/X _17173_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12048_/B sky130_fd_sc_hd__mux2_1
X_16924_ _17265_/CLK _16924_/D vssd1 vssd1 vccd1 vccd1 _16924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_193_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18374_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16855_ _18124_/CLK _16855_/D vssd1 vssd1 vccd1 vccd1 _16855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_122_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16131_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _17650_/CLK _15806_/D vssd1 vssd1 vccd1 vccd1 _15806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ _18019_/CLK _16786_/D vssd1 vssd1 vccd1 vccd1 _16786_/Q sky130_fd_sc_hd__dfxtp_1
X_13998_ _14894_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15737_ _17740_/CLK _15737_/D vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ hold3108/X hold3253/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _18456_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15668_ _17160_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17407_ _18456_/CLK _17407_/D vssd1 vssd1 vccd1 vccd1 _17407_/Q sky130_fd_sc_hd__dfxtp_1
X_14619_ hold2830/X _14612_/B _14618_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18387_ _18387_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15599_ _17215_/CLK _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08140_ hold181/A _15709_/Q hold240/A vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17338_ _17343_/CLK hold33/X vssd1 vssd1 vccd1 vccd1 _17338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ hold2976/X _08097_/A2 _08070_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _08071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _17269_/CLK _17269_/D vssd1 vssd1 vccd1 vccd1 _17269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4005 _15253_/X vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4016 _16369_/Q vssd1 vssd1 vccd1 vccd1 hold4016/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4027 _09790_/X vssd1 vssd1 vccd1 vccd1 _16420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4038 _17002_/Q vssd1 vssd1 vccd1 vccd1 hold4038/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3304 _17461_/Q vssd1 vssd1 vccd1 vccd1 hold3304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4049 _11359_/X vssd1 vssd1 vccd1 vccd1 _16943_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3315 _17482_/Q vssd1 vssd1 vccd1 vccd1 hold3315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3326 _16656_/Q vssd1 vssd1 vccd1 vccd1 hold3326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3337 _17442_/Q vssd1 vssd1 vccd1 vccd1 hold3337/X sky130_fd_sc_hd__dlygate4sd3_1
X_08973_ hold402/X hold480/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__mux2_1
Xhold2603 _16186_/Q vssd1 vssd1 vccd1 vccd1 hold2603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3348 _17436_/Q vssd1 vssd1 vccd1 vccd1 hold3348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3359 _16403_/Q vssd1 vssd1 vccd1 vccd1 hold3359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2614 _16270_/Q vssd1 vssd1 vccd1 vccd1 hold2614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__buf_4
XFILLER_0_209_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2625 _14203_/X vssd1 vssd1 vccd1 vccd1 _17902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2636 _17921_/Q vssd1 vssd1 vccd1 vccd1 hold2636/X sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _15547_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07924_/Y sky130_fd_sc_hd__nand2_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1902 _14454_/X vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 _17993_/Q vssd1 vssd1 vccd1 vccd1 hold2647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _14687_/X vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _15584_/Q vssd1 vssd1 vccd1 vccd1 hold2658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1924 _14895_/X vssd1 vssd1 vccd1 vccd1 _18234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 _15576_/Q vssd1 vssd1 vccd1 vccd1 hold2669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 _18185_/Q vssd1 vssd1 vccd1 vccd1 hold1935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1946 _14751_/X vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _15533_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__or2_1
Xhold1957 _14589_/X vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _18044_/Q vssd1 vssd1 vccd1 vccd1 hold1968/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1979 _15784_/Q vssd1 vssd1 vccd1 vccd1 hold1979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07786_ _07786_/A vssd1 vssd1 vccd1 vccd1 _07786_/Y sky130_fd_sc_hd__inv_2
X_09525_ _09987_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09463_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_0_231_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08407_ _15521_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08407_/X sky130_fd_sc_hd__or2_1
X_09387_ _15480_/A _09386_/X _18458_/Q vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08338_ hold764/A hold732/A hold329/X vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__or3_1
XFILLER_0_227_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08269_ hold2389/X _08268_/B _08268_/Y _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ hold5373/X _10625_/B _10299_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ _11694_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11280_/X sky130_fd_sc_hd__or2_1
Xhold5240 _16654_/Q vssd1 vssd1 vccd1 vccd1 hold5240/X sky130_fd_sc_hd__dlygate4sd3_1
X_10231_ hold5060/X _10637_/B _10230_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _10231_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5251 _11356_/X vssd1 vssd1 vccd1 vccd1 _16942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5262 _16686_/Q vssd1 vssd1 vccd1 vccd1 hold5262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5273 _12130_/X vssd1 vssd1 vccd1 vccd1 _17200_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5284 _16943_/Q vssd1 vssd1 vccd1 vccd1 hold5284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4550 _11608_/X vssd1 vssd1 vccd1 vccd1 _17026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5295 _11557_/X vssd1 vssd1 vccd1 vccd1 _17009_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10162_ hold3962/X _10622_/B _10161_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10162_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4561 _17712_/Q vssd1 vssd1 vccd1 vccd1 hold4561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4572 _15353_/X vssd1 vssd1 vccd1 vccd1 _15354_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4583 _17612_/Q vssd1 vssd1 vccd1 vccd1 hold4583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4594 _15453_/X vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3860 _16360_/Q vssd1 vssd1 vccd1 vccd1 hold3860/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ hold3659/X _10571_/B _10092_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10093_/X
+ sky130_fd_sc_hd__o211a_1
X_14970_ _15185_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__or2_1
Xhold3871 _11632_/X vssd1 vssd1 vccd1 vccd1 _17034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3882 _16649_/Q vssd1 vssd1 vccd1 vccd1 hold3882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3893 _10165_/X vssd1 vssd1 vccd1 vccd1 _16545_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _13921_/A _13921_/B vssd1 vssd1 vccd1 vccd1 _17766_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16640_ _18228_/CLK _16640_/D vssd1 vssd1 vccd1 vccd1 _16640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13852_ _13888_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _17737_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_230_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ hold3217/X _12802_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__mux2_1
X_16571_ _18223_/CLK _16571_/D vssd1 vssd1 vccd1 vccd1 _16571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13783_ hold4497/X _13877_/B _13782_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _13783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10995_ _11103_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10995_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18310_ _18349_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 hold471/A sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ hold2136/X _15560_/A2 _15521_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _15522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ hold3212/X _12733_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12735_/B sky130_fd_sc_hd__mux2_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ _18273_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15481_/A1 _15445_/X _15452_/X _15481_/B1 hold5876/A vssd1 vssd1 vccd1 vccd1
+ _15453_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_128_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ hold3800/X _12664_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14404_ hold2094/X _14446_/A2 _14403_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14404_/X
+ sky130_fd_sc_hd__o211a_1
X_18172_ _18210_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
X_11616_ _11712_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__or2_1
X_15384_ _15394_/A _15384_/B vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12596_ hold3233/X _12595_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ _17283_/CLK _17123_/D vssd1 vssd1 vccd1 vccd1 _17123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ hold2449/X _14326_/B _14334_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14335_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11547_ _11643_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__or2_1
Xhold509 hold509/A vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ _17900_/CLK _17054_/D vssd1 vssd1 vccd1 vccd1 _17054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14266_ _15541_/A _14266_/B vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11478_ _11670_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__or2_1
X_16005_ _18410_/CLK _16005_/D vssd1 vssd1 vccd1 vccd1 hold668/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13217_ _13217_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__and2_1
XFILLER_0_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10429_ hold5202/X _10619_/B _10428_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14197_ hold2160/X _14198_/B _14196_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _14197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_374_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17732_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ hold3591/X _13147_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__mux2_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_209_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13079_ _13199_/A1 _13077_/X _13078_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13079_/X
+ sky130_fd_sc_hd__o211a_2
X_17956_ _17996_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1209 _14017_/X vssd1 vssd1 vccd1 vccd1 _17812_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16907_ _18425_/CLK _16907_/D vssd1 vssd1 vccd1 vccd1 _16907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17887_ _17887_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16838_ _18039_/CLK _16838_/D vssd1 vssd1 vccd1 vccd1 _16838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16769_ _18068_/CLK _16769_/D vssd1 vssd1 vccd1 vccd1 _16769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ hold2488/X _09325_/B _09309_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _09310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09241_ _15517_/A hold2179/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18439_ _18452_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ _15555_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08123_ _08133_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_6_22_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_22_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08054_ _15513_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3101 _09304_/X vssd1 vssd1 vccd1 vccd1 _16262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3112 _18002_/Q vssd1 vssd1 vccd1 vccd1 hold3112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3123 _14753_/X vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3134 _18355_/Q vssd1 vssd1 vccd1 vccd1 hold3134/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2400 _07919_/X vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 _17471_/Q vssd1 vssd1 vccd1 vccd1 hold3145/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3156 _12539_/X vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 _15650_/Q vssd1 vssd1 vccd1 vccd1 hold2411/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2422 _15598_/Q vssd1 vssd1 vccd1 vccd1 hold2422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 _17477_/Q vssd1 vssd1 vccd1 vccd1 hold3167/X sky130_fd_sc_hd__dlygate4sd3_1
X_08956_ _12418_/A _08956_/B vssd1 vssd1 vccd1 vccd1 _16095_/D sky130_fd_sc_hd__and2_1
XFILLER_0_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3178 _12794_/X vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2433 _14273_/X vssd1 vssd1 vccd1 vccd1 _17935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2444 _14853_/X vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3189 _18088_/Q vssd1 vssd1 vccd1 vccd1 hold3189/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1710 _18221_/Q vssd1 vssd1 vccd1 vccd1 hold1710/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2455 _16160_/Q vssd1 vssd1 vccd1 vccd1 hold2455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2466 _14759_/X vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1721 _14277_/X vssd1 vssd1 vccd1 vccd1 _17937_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ hold2605/X _07924_/B _07906_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _07907_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1732 _14683_/X vssd1 vssd1 vccd1 vccd1 _18131_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2477 _17961_/Q vssd1 vssd1 vccd1 vccd1 hold2477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08887_ _15414_/A hold175/X vssd1 vssd1 vccd1 vccd1 _16061_/D sky130_fd_sc_hd__and2_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1743 _08259_/X vssd1 vssd1 vccd1 vccd1 _15764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2488 _16265_/Q vssd1 vssd1 vccd1 vccd1 hold2488/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2499 _14651_/X vssd1 vssd1 vccd1 vccd1 _18116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _14291_/X vssd1 vssd1 vccd1 vccd1 _17943_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1765 _18144_/Q vssd1 vssd1 vccd1 vccd1 hold1765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1776 _09095_/X vssd1 vssd1 vccd1 vccd1 _16162_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07838_ hold2729/X _07865_/B _07837_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07838_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1787 _18320_/Q vssd1 vssd1 vccd1 vccd1 hold1787/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1798 _14601_/X vssd1 vssd1 vccd1 vccd1 _18092_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ hold3968/X _10004_/B _09507_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09508_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ hold5585/X _11201_/B _10779_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _10780_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_6_61_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_61_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ hold1833/X _07804_/A _15304_/A _09438_/X vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _17318_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ hold5417/X _12329_/B _11400_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _11401_/X
+ sky130_fd_sc_hd__o211a_1
X_12381_ hold554/X hold704/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold705/A sky130_fd_sc_hd__mux2_1
XANTENNA_80 _17523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_91 hold746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _14854_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__or2_1
X_11332_ hold3762/X _11617_/A2 _11331_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14051_ hold1361/X _14038_/B _14050_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14051_/X
+ sky130_fd_sc_hd__o211a_1
X_11263_ hold5284/X _11747_/B _11262_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5070 _16677_/Q vssd1 vssd1 vccd1 vccd1 hold5070/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _17510_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5081 _13333_/X vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10214_ hold1927/X _16562_/Q _10580_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__mux2_1
Xhold5092 _16647_/Q vssd1 vssd1 vccd1 vccd1 hold5092/X sky130_fd_sc_hd__dlygate4sd3_1
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _16888_/D sky130_fd_sc_hd__nor2_1
XTAP_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4380 _16830_/Q vssd1 vssd1 vccd1 vccd1 hold4380/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ hold2971/X _16539_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4391 _17705_/Q vssd1 vssd1 vccd1 vccd1 hold4391/X sky130_fd_sc_hd__dlygate4sd3_1
X_17810_ _18426_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3690 _10099_/X vssd1 vssd1 vccd1 vccd1 _16523_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _17741_/CLK _17741_/D vssd1 vssd1 vccd1 vccd1 _17741_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ hold1117/X _14952_/B _14952_/Y _15028_/A vssd1 vssd1 vccd1 vccd1 _14953_/X
+ sky130_fd_sc_hd__o211a_1
X_10076_ hold1218/X hold3695/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_238_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _14854_/A hold1348/X hold124/X vssd1 vssd1 vccd1 vccd1 _13905_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_215_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17672_ _17736_/CLK _17672_/D vssd1 vssd1 vccd1 vccd1 _17672_/Q sky130_fd_sc_hd__dfxtp_1
X_14884_ hold972/X _14894_/B vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16623_ _18153_/CLK _16623_/D vssd1 vssd1 vccd1 vccd1 _16623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _17732_/Q _13856_/B _13856_/C vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__and3_1
XFILLER_0_98_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16554_ _18142_/CLK _16554_/D vssd1 vssd1 vccd1 vccd1 _16554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ hold2791/X hold5691/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ hold5551/X _11732_/B _10977_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _10978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ _15521_/A hold1987/X hold691/X vssd1 vssd1 vccd1 vccd1 _15506_/B sky130_fd_sc_hd__mux2_1
X_12717_ _12759_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _17415_/D sky130_fd_sc_hd__and2_1
X_16485_ _18300_/CLK _16485_/D vssd1 vssd1 vccd1 vccd1 _16485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ hold2000/X hold5214/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13698_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _18224_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15436_ _17319_/Q _09357_/A _09392_/A hold758/X vssd1 vssd1 vccd1 vccd1 _15436_/X
+ sky130_fd_sc_hd__a22o_1
X_12648_ _12654_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _17392_/D sky130_fd_sc_hd__and2_1
X_18155_ _18219_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15367_ _16145_/Q _15487_/A2 _15484_/B1 hold128/X _15366_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_182_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _12969_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _17369_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _17266_/CLK _17106_/D vssd1 vssd1 vccd1 vccd1 _17106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _15105_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _18234_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ _15943_/Q _15484_/A2 _09392_/D hold421/X vssd1 vssd1 vccd1 vccd1 _15298_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold328 hold688/X vssd1 vssd1 vccd1 vccd1 hold689/A sky130_fd_sc_hd__buf_4
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _17883_/CLK _17037_/D vssd1 vssd1 vccd1 vccd1 _17037_/Q sky130_fd_sc_hd__dfxtp_1
X_14249_ hold1632/X _14266_/B _14248_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout808 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _14829_/C1 sky130_fd_sc_hd__buf_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__buf_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ hold113/X _16024_/Q _08866_/S vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__mux2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ hold4026/X _11201_/B _09789_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09790_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _15823_/Q vssd1 vssd1 vccd1 vccd1 hold1006/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _08366_/X vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ hold17/X hold477/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__mux2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 hold1033/X vssd1 vssd1 vccd1 vccd1 hold1034/A sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ _17971_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1039 _14227_/X vssd1 vssd1 vccd1 vccd1 _17913_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08672_ _12426_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _15553_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ hold2923/X _09177_/A2 _09154_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08106_ hold999/X hold1023/X hold240/X vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_296_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17999_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ hold944/X _09098_/B vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_225_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18163_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08037_ _14330_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08037_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold840 hold840/A vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold851 hold851/A vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold884 hold884/A vssd1 vssd1 vccd1 vccd1 hold884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 hold895/A vssd1 vssd1 vccd1 vccd1 hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _13078_/A _10004_/B _09987_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09988_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2230 _08208_/X vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _14123_/X vssd1 vssd1 vccd1 vccd1 _17863_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2252 _18096_/Q vssd1 vssd1 vccd1 vccd1 hold2252/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08939_ hold215/X hold883/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold884/A sky130_fd_sc_hd__mux2_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2263 _14436_/X vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2274 _17861_/Q vssd1 vssd1 vccd1 vccd1 hold2274/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2285 _15170_/X vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1540 _15566_/Q vssd1 vssd1 vccd1 vccd1 hold1540/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1551 la_data_in[14] vssd1 vssd1 vccd1 vccd1 hold1551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2296 _08428_/X vssd1 vssd1 vccd1 vccd1 _15844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ hold4233/X _13868_/B _11949_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _11950_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1562 _14057_/X vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1573 _18361_/Q vssd1 vssd1 vccd1 vccd1 hold1573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1584 _09292_/X vssd1 vssd1 vccd1 vccd1 _16256_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ hold1701/X _16791_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__mux2_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1595 _15869_/Q vssd1 vssd1 vccd1 vccd1 hold1595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ hold4221/X _13871_/B _11880_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _13716_/A _13620_/B vssd1 vssd1 vccd1 vccd1 _13620_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ hold1397/X hold5192/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _13761_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__or2_1
X_10763_ hold1003/X hold3476/X _11147_/C vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _17344_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16270_ _17372_/CLK _16270_/D vssd1 vssd1 vccd1 vccd1 _16270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13482_ _13698_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13482_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ hold1632/X hold3691/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15221_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__nand2_1
X_12433_ hold210/X hold322/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__mux2_1
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15152_ hold6002/X _15167_/B hold1048/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__o211a_1
X_12364_ _13873_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _17278_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14103_ hold2763/X _14107_/A2 _14102_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _14103_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ hold2559/X hold3670/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__mux2_1
X_15083_ _15191_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ _13825_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _17255_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _15541_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nand2_1
X_11246_ hold1987/X hold3563/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11177_ _16883_/Q _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10128_ _10536_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10128_/X sky130_fd_sc_hd__or2_1
XTAP_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15985_ _17347_/CLK _15985_/D vssd1 vssd1 vccd1 vccd1 _15985_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10059_ _13270_/A _10191_/A _10058_/X vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__a21oi_1
X_14936_ _15205_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14936_/X sky130_fd_sc_hd__or2_1
X_17724_ _17724_/CLK _17724_/D vssd1 vssd1 vccd1 vccd1 _17724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17509_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14867_ hold1147/X _14882_/B _14866_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14867_/X
+ sky130_fd_sc_hd__o211a_1
X_17655_ _17693_/CLK _17655_/D vssd1 vssd1 vccd1 vccd1 _17655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _18182_/CLK _16606_/D vssd1 vssd1 vccd1 vccd1 _16606_/Q sky130_fd_sc_hd__dfxtp_1
X_13818_ hold4643/X _13698_/A _13817_/X vssd1 vssd1 vccd1 vccd1 _13818_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17586_ _17746_/CLK _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14798_ _15191_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__or2_1
XFILLER_0_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ _18163_/CLK _16537_/D vssd1 vssd1 vccd1 vccd1 _16537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13749_ _13788_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16468_ _18379_/CLK _16468_/D vssd1 vssd1 vccd1 vccd1 _16468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18207_ _18262_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
X_15419_ hold413/X _09386_/A _15417_/X vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16399_ _18342_/CLK _16399_/D vssd1 vssd1 vccd1 vccd1 _16399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18138_ _18170_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5806 hold5806/A vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_12
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5817 _18405_/Q vssd1 vssd1 vccd1 vccd1 hold5817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 hold243/X vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5828 _17518_/Q vssd1 vssd1 vccd1 vccd1 hold990/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5839 _17520_/Q vssd1 vssd1 vccd1 vccd1 hold5839/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18069_ _18071_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ hold1811/X hold3802/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__mux2_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout605 _09364_/Y vssd1 vssd1 vccd1 vccd1 _15451_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout616 _09354_/Y vssd1 vssd1 vccd1 vccd1 _15487_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ hold3139/X _16438_/Q _10034_/C vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout627 hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout638 _12696_/A vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout649 _12804_/A vssd1 vssd1 vccd1 vccd1 _15548_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_225_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09773_ hold1074/X hold3613/X _10601_/C vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__mux2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _09053_/A hold299/X vssd1 vssd1 vccd1 vccd1 _15983_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ hold140/X hold286/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08586_ hold145/X hold158/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09207_ hold1216/X _09216_/B _09206_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _09207_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_406_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17883_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09138_ _15521_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ hold6000/X _09119_/A2 hold1113/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ hold1684/X _17184_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__mux2_1
Xhold670 hold670/A vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 hold743/X vssd1 vssd1 vccd1 vccd1 hold744/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold692 hold692/A vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _11124_/A _11031_/B vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 _17773_/Q vssd1 vssd1 vccd1 vccd1 hold2060/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _08308_/X vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15770_ _17689_/CLK _15770_/D vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2082 _15518_/X vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ hold2184/X hold3136/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__mux2_1
Xhold2093 _14329_/X vssd1 vssd1 vccd1 vccd1 _17962_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 _07989_/X vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 _16287_/Q vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__buf_1
X_14721_ hold2492/X _14720_/B _14720_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14721_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ hold2976/X _17135_/Q _12314_/C vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__mux2_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _14099_/X vssd1 vssd1 vccd1 vccd1 _17852_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _18435_/CLK _17440_/D vssd1 vssd1 vccd1 vccd1 _17440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _15099_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14652_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11864_ hold1609/X hold3825/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__mux2_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ hold5214/X _13817_/B _13602_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13603_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17372_/CLK _17371_/D vssd1 vssd1 vccd1 vccd1 _17371_/Q sky130_fd_sc_hd__dfxtp_1
X_10815_ _11124_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__or2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ hold2291/X _14610_/B _14582_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11795_ _17089_/Q _12365_/B _12365_/C vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__and3_1
XFILLER_0_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16322_ _16322_/CLK _16322_/D vssd1 vssd1 vccd1 vccd1 hold895/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13534_ hold5707/X _13829_/B _13533_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13534_/X
+ sky130_fd_sc_hd__o211a_1
X_10746_ _11670_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_147_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18373_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16253_ _17435_/CLK _16253_/D vssd1 vssd1 vccd1 vccd1 _16253_/Q sky130_fd_sc_hd__dfxtp_1
X_13465_ hold4521/X _13777_/A2 _13464_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10677_ _11064_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15204_ hold1648/X _15221_/B _15203_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _15204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12416_ _12416_/A _12416_/B vssd1 vssd1 vccd1 vccd1 _17301_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16184_ _17469_/CLK _16184_/D vssd1 vssd1 vccd1 vccd1 _16184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13396_ hold4389/X _13886_/B _13395_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15135_ _15189_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ _12347_/A _12347_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _15066_/A _15066_/B vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12278_ hold1239/X hold4151/X _13556_/S vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ hold1208/X _14040_/B _14016_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _14017_/X
+ sky130_fd_sc_hd__o211a_1
X_11229_ _12213_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _18401_/CLK _15968_/D vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17707_ _17707_/CLK _17707_/D vssd1 vssd1 vccd1 vccd1 _17707_/Q sky130_fd_sc_hd__dfxtp_1
X_14919_ hold1799/X _14946_/B _14918_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14919_/X
+ sky130_fd_sc_hd__o211a_1
X_15899_ _17303_/CLK _15899_/D vssd1 vssd1 vccd1 vccd1 hold706/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08440_ hold2482/X _08440_/A2 _08439_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17638_ _17702_/CLK _17638_/D vssd1 vssd1 vccd1 vccd1 _17638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08379_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _15817_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17569_ _17728_/CLK _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5603 _16992_/Q vssd1 vssd1 vccd1 vccd1 hold5603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5614 _11695_/X vssd1 vssd1 vccd1 vccd1 _17055_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5625 _16827_/Q vssd1 vssd1 vccd1 vccd1 hold5625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5636 _11011_/X vssd1 vssd1 vccd1 vccd1 _16827_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4902 _10090_/X vssd1 vssd1 vccd1 vccd1 _16520_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5647 _17015_/Q vssd1 vssd1 vccd1 vccd1 hold5647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5658 _13830_/Y vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4913 _17223_/Q vssd1 vssd1 vccd1 vccd1 hold4913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4924 _10555_/X vssd1 vssd1 vccd1 vccd1 _16675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5669 _16382_/Q vssd1 vssd1 vccd1 vccd1 hold5669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4935 _13435_/X vssd1 vssd1 vccd1 vccd1 _17598_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4946 _17252_/Q vssd1 vssd1 vccd1 vccd1 hold4946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4957 _12202_/X vssd1 vssd1 vccd1 vccd1 _17224_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4968 _16653_/Q vssd1 vssd1 vccd1 vccd1 hold4968/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout402 hold332/X vssd1 vssd1 vccd1 vccd1 _14391_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_239_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4979 _10363_/X vssd1 vssd1 vccd1 vccd1 _16611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout413 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__buf_8
Xfanout424 hold123/X vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__buf_6
Xfanout435 _12302_/C vssd1 vssd1 vccd1 vccd1 _13412_/S sky130_fd_sc_hd__buf_6
Xfanout446 _11711_/S vssd1 vssd1 vccd1 vccd1 _12308_/C sky130_fd_sc_hd__buf_6
X_09825_ _09843_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__or2_1
Xfanout457 _13847_/C vssd1 vssd1 vccd1 vccd1 _13856_/C sky130_fd_sc_hd__buf_6
Xfanout468 _12368_/C vssd1 vssd1 vccd1 vccd1 _13877_/C sky130_fd_sc_hd__buf_6
Xfanout479 _11219_/C vssd1 vssd1 vccd1 vccd1 _11768_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09756_ _09936_/A _09756_/B vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08707_ hold228/X hold702/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__mux2_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09687_ _10191_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__or2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _12416_/A hold540/X vssd1 vssd1 vccd1 vccd1 _15941_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08569_ _09055_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _15908_/D sky130_fd_sc_hd__and2_1
XFILLER_0_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ _11194_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _16690_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _12243_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10531_ hold4863/X _10625_/B _10530_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_240_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18152_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _17582_/Q _17116_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__mux2_1
X_10462_ hold3643/X _11180_/B _10461_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ _13716_/A _12201_/B vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__or2_1
X_13181_ _13180_/X hold4636/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ hold4968/X _10601_/B _10392_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ _12267_/A _12132_/B vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12063_ _12231_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or2_1
X_16940_ _17822_/CLK _16940_/D vssd1 vssd1 vccd1 vccd1 _16940_/Q sky130_fd_sc_hd__dfxtp_1
X_11014_ hold4427/X _11210_/B _11013_/X _14538_/C1 vssd1 vssd1 vccd1 vccd1 _11014_/X
+ sky130_fd_sc_hd__o211a_1
X_16871_ _18042_/CLK _16871_/D vssd1 vssd1 vccd1 vccd1 _16871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _17701_/CLK _15822_/D vssd1 vssd1 vccd1 vccd1 _15822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _17736_/CLK _15753_/D vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ hold3289/X _12964_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__mux2_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14704_ _14758_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__or2_1
X_11916_ _12204_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_399_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17834_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_213_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15684_ _17872_/CLK _15684_/D vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12896_ hold3377/X _12895_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__mux2_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14635_ hold2941/X _14666_/B _14634_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _14635_/X
+ sky130_fd_sc_hd__o211a_1
X_17423_ _17689_/CLK _17423_/D vssd1 vssd1 vccd1 vccd1 _17423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_328_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17808_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ _12267_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__or2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ hold690/X _14573_/B hold2006/X vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__a21o_1
X_17354_ _17378_/CLK _17354_/D vssd1 vssd1 vccd1 vccd1 _17354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ hold4689/X _12285_/A _11777_/X vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16305_ _18404_/CLK _16305_/D vssd1 vssd1 vccd1 vccd1 _16305_/Q sky130_fd_sc_hd__dfxtp_1
X_13517_ _15811_/Q hold4010/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__mux2_1
X_17285_ _17301_/CLK _17285_/D vssd1 vssd1 vccd1 vccd1 hold340/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10729_ hold4509/X _11768_/B _10728_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14497_ _15231_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16236_ _17429_/CLK _16236_/D vssd1 vssd1 vccd1 vccd1 _16236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ hold2869/X hold5735/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16167_ _17879_/CLK _16167_/D vssd1 vssd1 vccd1 vccd1 _16167_/Q sky130_fd_sc_hd__dfxtp_1
X_13379_ hold1595/X hold3649/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__mux2_1
Xhold4209 _17721_/Q vssd1 vssd1 vccd1 vccd1 hold4209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15118_ hold5993/X _15113_/B hold560/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 hold561/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16098_ _16126_/CLK _16098_/D vssd1 vssd1 vccd1 vccd1 hold811/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3508 _17419_/Q vssd1 vssd1 vccd1 vccd1 hold3508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3519 _17685_/Q vssd1 vssd1 vccd1 vccd1 hold3519/X sky130_fd_sc_hd__dlygate4sd3_1
X_15049_ _15103_/A hold3038/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__mux2_1
X_07940_ _14164_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__or2_1
XFILLER_0_220_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2807 _09151_/X vssd1 vssd1 vccd1 vccd1 _16188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2818 _17974_/Q vssd1 vssd1 vccd1 vccd1 hold2818/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2829 _07945_/X vssd1 vssd1 vccd1 vccd1 _15615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17875_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07871_ _15549_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07871_/X sky130_fd_sc_hd__or2_1
X_09610_ hold3966/X _10004_/B _09609_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09610_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09541_ hold4016/X _10019_/B _09540_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09541_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09472_ _09472_/A _09472_/B _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09477_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_149_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _15211_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08423_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08354_ _15523_/A _15809_/Q hold134/X vssd1 vssd1 vccd1 vccd1 _08354_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08285_ _14164_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5400 _09622_/X vssd1 vssd1 vccd1 vccd1 _16364_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5411 _16941_/Q vssd1 vssd1 vccd1 vccd1 hold5411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5422 _12262_/X vssd1 vssd1 vccd1 vccd1 _17244_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5433 _16569_/Q vssd1 vssd1 vccd1 vccd1 hold5433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5444 _11878_/X vssd1 vssd1 vccd1 vccd1 _17116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4710 _09775_/X vssd1 vssd1 vccd1 vccd1 _16415_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5455 _17243_/Q vssd1 vssd1 vccd1 vccd1 hold5455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4721 _16684_/Q vssd1 vssd1 vccd1 vccd1 hold4721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5466 _11974_/X vssd1 vssd1 vccd1 vccd1 _17148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4732 _09586_/X vssd1 vssd1 vccd1 vccd1 _16352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5477 _16772_/Q vssd1 vssd1 vccd1 vccd1 hold5477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4743 _16404_/Q vssd1 vssd1 vccd1 vccd1 hold4743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5488 _10849_/X vssd1 vssd1 vccd1 vccd1 _16773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4754 _10798_/X vssd1 vssd1 vccd1 vccd1 _16756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5499 _17613_/Q vssd1 vssd1 vccd1 vccd1 hold5499/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4765 _16448_/Q vssd1 vssd1 vccd1 vccd1 hold4765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4776 _10081_/X vssd1 vssd1 vccd1 vccd1 _16517_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout210 _10019_/B vssd1 vssd1 vccd1 vccd1 _11156_/B sky130_fd_sc_hd__buf_4
Xfanout221 _11192_/B vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__buf_4
Xhold4787 _17101_/Q vssd1 vssd1 vccd1 vccd1 hold4787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4798 _09961_/X vssd1 vssd1 vccd1 vccd1 _16477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout232 fanout246/X vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__buf_4
XFILLER_0_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout243 _10637_/B vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__clkbuf_8
Xfanout254 _13623_/A vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__buf_4
Xfanout265 _11652_/A vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__buf_4
XFILLER_0_195_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout276 fanout334/X vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__buf_4
X_09808_ hold5110/X _11159_/B _09807_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09808_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout287 _12051_/A vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__clkbuf_4
Xfanout298 _09843_/A vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__buf_4
XFILLER_0_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ hold3386/X _10007_/B _09738_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09739_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12750_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _17426_/D sky130_fd_sc_hd__and2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11701_ hold4327/X _12365_/B _11700_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11701_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_421_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12780_/A _12681_/B vssd1 vssd1 vccd1 vccd1 _17403_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ hold3041/X _14433_/B _14419_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _14420_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ hold3870/X _11726_/B _11631_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ hold525/A _17973_/Q hold333/X vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__mux2_1
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ hold5529/X _11753_/B _11562_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _13302_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ hold2546/X _16662_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__mux2_1
X_17070_ _17852_/CLK _17070_/D vssd1 vssd1 vccd1 vccd1 _17070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14282_ _14443_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__or2_1
X_11494_ hold5124/X _12314_/B _11493_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11494_/X
+ sky130_fd_sc_hd__o211a_1
X_16021_ _17313_/CLK _16021_/D vssd1 vssd1 vccd1 vccd1 hold773/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13233_ _13233_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__and2_1
XFILLER_0_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10445_ hold2935/X hold4974/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ hold4660/X _13163_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__mux2_2
X_10376_ hold1921/X hold4757/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12115_ hold5096/X _12308_/B _12114_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _12115_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13095_ _13199_/A1 _13093_/X _13094_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13095_/X
+ sky130_fd_sc_hd__o211a_1
X_17972_ _18035_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
X_12046_ hold4235/X _13868_/B _12045_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__o211a_1
X_16923_ _17769_/CLK _16923_/D vssd1 vssd1 vccd1 vccd1 _16923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16854_ _18055_/CLK _16854_/D vssd1 vssd1 vccd1 vccd1 _16854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _17642_/CLK _15805_/D vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfxtp_1
X_13997_ hold1287/X _13986_/B _13996_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13997_/X
+ sky130_fd_sc_hd__o211a_1
X_16785_ _18018_/CLK _16785_/D vssd1 vssd1 vccd1 vccd1 _16785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _12990_/A _12948_/B vssd1 vssd1 vccd1 vccd1 _17492_/D sky130_fd_sc_hd__and2_1
X_15736_ _17701_/CLK _15736_/D vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_162_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18309_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_213_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18455_ _18455_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
X_15667_ _17221_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12990_/A _12879_/B vssd1 vssd1 vccd1 vccd1 _17469_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17406_ _18455_/CLK _17406_/D vssd1 vssd1 vccd1 vccd1 _17406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14618_ _14726_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__or2_1
X_18386_ _18386_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _17234_/CLK _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17337_ _17339_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 _17337_/Q sky130_fd_sc_hd__dfxtp_1
X_14549_ _15229_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_12_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_12_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _15529_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ _17711_/CLK _17268_/D vssd1 vssd1 vccd1 vccd1 _17268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ _17481_/CLK _16219_/D vssd1 vssd1 vccd1 vccd1 _16219_/Q sky130_fd_sc_hd__dfxtp_1
X_17199_ _17199_/CLK _17199_/D vssd1 vssd1 vccd1 vccd1 _17199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4006 _16431_/Q vssd1 vssd1 vccd1 vccd1 hold4006/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4017 _09541_/X vssd1 vssd1 vccd1 vccd1 _16337_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4028 _16645_/Q vssd1 vssd1 vccd1 vccd1 hold4028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4039 _11440_/X vssd1 vssd1 vccd1 vccd1 _16970_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3305 _12854_/X vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3316 _12917_/X vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _09055_/A _08972_/B vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__and2_1
Xhold3327 _10402_/X vssd1 vssd1 vccd1 vccd1 _16624_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3338 _17435_/Q vssd1 vssd1 vccd1 vccd1 hold3338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3349 _16457_/Q vssd1 vssd1 vccd1 vccd1 hold3349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2604 _09147_/X vssd1 vssd1 vccd1 vccd1 _16186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 _09320_/X vssd1 vssd1 vccd1 vccd1 _16270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ hold2441/X _07924_/B _07922_/Y _08163_/A vssd1 vssd1 vccd1 vccd1 _07923_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2626 _16194_/Q vssd1 vssd1 vccd1 vccd1 hold2626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2637 _14245_/X vssd1 vssd1 vccd1 vccd1 _17921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 _17981_/Q vssd1 vssd1 vccd1 vccd1 hold1903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _15654_/Q vssd1 vssd1 vccd1 vccd1 hold2648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 _18224_/Q vssd1 vssd1 vccd1 vccd1 hold1914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _07878_/X vssd1 vssd1 vccd1 vccd1 _15584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 _17823_/Q vssd1 vssd1 vccd1 vccd1 hold1925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1936 _14795_/X vssd1 vssd1 vccd1 vccd1 _18185_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07854_ hold2286/X _07869_/B _07853_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07854_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1947 _18456_/Q vssd1 vssd1 vccd1 vccd1 hold1947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1958 _17942_/Q vssd1 vssd1 vccd1 vccd1 hold1958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 _14498_/X vssd1 vssd1 vccd1 vccd1 _18044_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07785_ _09438_/B vssd1 vssd1 vccd1 vccd1 _07785_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ hold1591/X _13126_/A _10004_/C vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_6_51_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_51_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09456_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09457_/C sky130_fd_sc_hd__or2_1
XFILLER_0_148_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ hold1225/X _08440_/A2 _08405_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08406_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09386_ _09386_/A _09386_/B _09392_/C _09386_/D vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_164_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08337_ hold752/A hold689/A vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__nand2_1
XFILLER_0_191_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08268_ _15547_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08199_ _15533_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5230 _17052_/Q vssd1 vssd1 vccd1 vccd1 hold5230/X sky130_fd_sc_hd__dlygate4sd3_1
X_10230_ _10542_/A _10230_/B vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__or2_1
Xhold5241 _10396_/X vssd1 vssd1 vccd1 vccd1 _16622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5252 _16490_/Q vssd1 vssd1 vccd1 vccd1 hold5252/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5263 _10492_/X vssd1 vssd1 vccd1 vccd1 _16654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5274 _17222_/Q vssd1 vssd1 vccd1 vccd1 hold5274/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4540 _10933_/X vssd1 vssd1 vccd1 vccd1 _16801_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5285 _11263_/X vssd1 vssd1 vccd1 vccd1 _16911_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10161_ _10527_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10161_/X sky130_fd_sc_hd__or2_1
Xhold5296 _17262_/Q vssd1 vssd1 vccd1 vccd1 hold5296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4551 _17208_/Q vssd1 vssd1 vccd1 vccd1 hold4551/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4562 _13681_/X vssd1 vssd1 vccd1 vccd1 _17680_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4573 hold5887/X vssd1 vssd1 vccd1 vccd1 hold5888/A sky130_fd_sc_hd__buf_6
XFILLER_0_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4584 _13381_/X vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4595 _16343_/Q vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3850 _16737_/Q vssd1 vssd1 vccd1 vccd1 hold3850/X sky130_fd_sc_hd__buf_1
Xhold3861 _09514_/X vssd1 vssd1 vccd1 vccd1 _16328_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10092_ _10470_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3872 _16664_/Q vssd1 vssd1 vccd1 vccd1 hold3872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3883 _10381_/X vssd1 vssd1 vccd1 vccd1 _16617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3894 _16778_/Q vssd1 vssd1 vccd1 vccd1 hold3894/X sky130_fd_sc_hd__dlygate4sd3_1
X_13920_ _14529_/A hold1349/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__mux2_1
X_13851_ hold3697/X _13791_/A _13850_/X vssd1 vssd1 vccd1 vccd1 _13851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_236_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12802_ hold2242/X _17445_/Q _12826_/S vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16570_ _18222_/CLK _16570_/D vssd1 vssd1 vccd1 vccd1 _16570_/Q sky130_fd_sc_hd__dfxtp_1
X_13782_ _13782_/A _13782_/B vssd1 vssd1 vccd1 vccd1 _13782_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ hold3234/X _16822_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ hold2663/X hold3211/X _12748_/S vssd1 vssd1 vccd1 vccd1 _12733_/X sky130_fd_sc_hd__mux2_1
X_15521_ _15521_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _15489_/A _15452_/B _15452_/C _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/X
+ sky130_fd_sc_hd__or4_1
X_18240_ _18413_/CLK hold527/X vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ hold2040/X hold3770/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__mux2_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14403_ _14403_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ hold2540/X hold3746/X _11711_/S vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18171_ _18205_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
X_15383_ _15481_/A1 _15375_/X _15382_/X _15490_/B1 hold5848/A vssd1 vssd1 vccd1 vccd1
+ _15383_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ hold2418/X hold3227/X _12967_/S vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17122_ _17237_/CLK _17122_/D vssd1 vssd1 vccd1 vccd1 _17122_/Q sky130_fd_sc_hd__dfxtp_1
X_14334_ _14782_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14334_/X sky130_fd_sc_hd__or2_1
X_11546_ hold1391/X hold5222/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17053_ _17804_/CLK _17053_/D vssd1 vssd1 vccd1 vccd1 _17053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ hold2842/X _14272_/B _14264_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14265_/X
+ sky130_fd_sc_hd__o211a_1
X_11477_ hold1361/X hold5637/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ _18409_/CLK _16004_/D vssd1 vssd1 vccd1 vccd1 _16004_/Q sky130_fd_sc_hd__dfxtp_1
X_13216_ _13209_/X _13215_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17545_/D sky130_fd_sc_hd__o21a_1
X_10428_ _10524_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14196_ _14946_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13146_/X hold5917/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ _10527_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ _13078_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__or2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _18018_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12029_ hold2321/X _17167_/Q _12029_/S vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__mux2_1
X_16906_ _18430_/CLK _16906_/D vssd1 vssd1 vccd1 vccd1 _16906_/Q sky130_fd_sc_hd__dfxtp_1
X_17886_ _17886_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _18038_/CLK _16837_/D vssd1 vssd1 vccd1 vccd1 _16837_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_343_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17650_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_178_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16768_ _18065_/CLK _16768_/D vssd1 vssd1 vccd1 vccd1 _16768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15719_ _17719_/CLK _15719_/D vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16699_ _18223_/CLK _16699_/D vssd1 vssd1 vccd1 vccd1 _16699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09240_ _12768_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _16231_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438_ _18438_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09171_ hold2768/X _09177_/A2 _09170_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _18395_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08122_ _14862_/A hold2168/X hold240/X vssd1 vssd1 vccd1 vccd1 _08123_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08053_ hold1098/X _08097_/A2 _08052_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3102 _15621_/Q vssd1 vssd1 vccd1 vccd1 hold3102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3113 _14412_/X vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3124 _18003_/Q vssd1 vssd1 vccd1 vccd1 hold3124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3135 _15148_/X vssd1 vssd1 vccd1 vccd1 _18355_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2401 _16218_/Q vssd1 vssd1 vccd1 vccd1 hold2401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3146 _12884_/X vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08955_ hold98/X hold660/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__mux2_1
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3157 _17353_/Q vssd1 vssd1 vccd1 vccd1 hold3157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2412 _08018_/X vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 _18251_/Q vssd1 vssd1 vccd1 vccd1 hold3168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 _07909_/X vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3179 _17452_/Q vssd1 vssd1 vccd1 vccd1 hold3179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 _17847_/Q vssd1 vssd1 vccd1 vccd1 hold2434/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2445 _15753_/Q vssd1 vssd1 vccd1 vccd1 hold2445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 _13975_/X vssd1 vssd1 vccd1 vccd1 _17792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 _14869_/X vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _15529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__or2_1
Xhold2456 _09091_/X vssd1 vssd1 vccd1 vccd1 _16160_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08886_ hold174/X _16061_/Q _08928_/S vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__mux2_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1722 hold1889/X vssd1 vssd1 vccd1 vccd1 hold1890/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2467 _17840_/Q vssd1 vssd1 vccd1 vccd1 hold2467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _18353_/Q vssd1 vssd1 vccd1 vccd1 hold1733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _14327_/X vssd1 vssd1 vccd1 vccd1 _17961_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2489 _09310_/X vssd1 vssd1 vccd1 vccd1 _16265_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1744 _15879_/Q vssd1 vssd1 vccd1 vccd1 hold1744/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1755 _15801_/Q vssd1 vssd1 vccd1 vccd1 hold1755/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1766 _14709_/X vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07837_ _15515_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07837_/X sky130_fd_sc_hd__or2_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1777 _16315_/Q vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _15076_/X vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1799 _18244_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _09987_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09438_ _16305_/Q _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09369_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_240_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _12234_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12380_ _12380_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12401_/S sky130_fd_sc_hd__or2_2
XFILLER_0_35_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_70 hold998/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _15551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 hold746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11331_ _11712_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _14443_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14050_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _11652_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5060 _16599_/Q vssd1 vssd1 vccd1 vccd1 hold5060/X sky130_fd_sc_hd__dlygate4sd3_1
X_13001_ hold3609/X _13000_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__mux2_1
X_10213_ hold4925/X _10619_/B _10212_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5071 _10465_/X vssd1 vssd1 vccd1 vccd1 _16645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5082 _16600_/Q vssd1 vssd1 vccd1 vccd1 hold5082/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5093 _10375_/X vssd1 vssd1 vccd1 vccd1 _16615_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11193_ hold4625/X _11100_/A _11192_/X vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4370 _17248_/Q vssd1 vssd1 vccd1 vccd1 hold4370/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10144_ hold3789/X _10622_/B _10143_/X _14805_/C1 vssd1 vssd1 vccd1 vccd1 _10144_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4381 _10924_/X vssd1 vssd1 vccd1 vccd1 _16798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4392 _13660_/X vssd1 vssd1 vccd1 vccd1 _17673_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3680 _11145_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _17740_/CLK _17740_/D vssd1 vssd1 vccd1 vccd1 _17740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ _10603_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _16515_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_175_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _15221_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nand2_1
Xhold3691 _16722_/Q vssd1 vssd1 vccd1 vccd1 hold3691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2990 _14851_/X vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13903_ _13903_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _17757_/D sky130_fd_sc_hd__and2_1
X_17671_ _17703_/CLK _17671_/D vssd1 vssd1 vccd1 vccd1 _17671_/Q sky130_fd_sc_hd__dfxtp_1
X_14883_ hold1279/X _14882_/B _14882_/Y _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14883_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16622_ _18178_/CLK _16622_/D vssd1 vssd1 vccd1 vccd1 _16622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _13864_/A _13834_/B vssd1 vssd1 vccd1 vccd1 _17731_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_199_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _18141_/CLK _16553_/D vssd1 vssd1 vccd1 vccd1 _16553_/Q sky130_fd_sc_hd__dfxtp_1
X_13765_ hold4207/X _13883_/B _13764_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13765_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10977_ _11553_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ _15506_/A hold692/X vssd1 vssd1 vccd1 vccd1 hold693/A sky130_fd_sc_hd__and2_1
XFILLER_0_112_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12716_ hold3410/X _12715_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__mux2_1
X_16484_ _18395_/CLK _16484_/D vssd1 vssd1 vccd1 vccd1 _16484_/Q sky130_fd_sc_hd__dfxtp_1
X_13696_ hold4330/X _13886_/B _13695_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18223_ _18223_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ hold188/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ hold3799/X _12646_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ _17340_/Q _15448_/B1 _15485_/B1 _16117_/Q vssd1 vssd1 vccd1 vccd1 _15366_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18154_ _18154_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12578_ hold3170/X _12577_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17105_ _17265_/CLK _17105_/D vssd1 vssd1 vccd1 vccd1 _17105_/Q sky130_fd_sc_hd__dfxtp_1
X_14317_ hold3110/X hold756/X _14316_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14317_/X
+ sky130_fd_sc_hd__o211a_1
X_11529_ _12204_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__or2_1
X_15297_ hold544/X _15487_/A2 _15484_/B1 hold598/X _15296_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/B sky130_fd_sc_hd__a221o_1
X_18085_ _18113_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14248_ _14517_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14248_/X sky130_fd_sc_hd__or2_1
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ _17882_/CLK _17036_/D vssd1 vssd1 vccd1 vccd1 _17036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ hold1468/X _14202_/B _14178_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _14179_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 fanout847/X vssd1 vssd1 vccd1 vccd1 _09976_/C1 sky130_fd_sc_hd__buf_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _12444_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _15990_/D sky130_fd_sc_hd__and2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 hold1104/X vssd1 vssd1 vccd1 vccd1 hold1105/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 hold1045/X vssd1 vssd1 vccd1 vccd1 hold1046/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _18003_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1029 hold1035/X vssd1 vssd1 vccd1 vccd1 hold1029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08671_ hold113/X hold785/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17869_ _17869_/CLK _17869_/D vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ hold1375/X _09216_/B _09222_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09154_ _15537_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08105_ _15498_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _15691_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09085_ hold3108/X _09119_/A2 _09084_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09085_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08036_ hold2149/X _08033_/B _08035_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _08036_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold830 hold830/A vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold841 hold841/A vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold885 hold885/A vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold896 hold896/A vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_265_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18032_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__or2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2220 _15711_/Q vssd1 vssd1 vccd1 vccd1 hold2220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2231 _15874_/Q vssd1 vssd1 vccd1 vccd1 hold2231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _15324_/A hold550/X vssd1 vssd1 vccd1 vccd1 _16086_/D sky130_fd_sc_hd__and2_1
XFILLER_0_157_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2242 _16213_/Q vssd1 vssd1 vccd1 vccd1 hold2242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2253 _14609_/X vssd1 vssd1 vccd1 vccd1 _18096_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2264 _15824_/Q vssd1 vssd1 vccd1 vccd1 hold2264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1530 _14731_/X vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2275 _14119_/X vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1541 _07842_/X vssd1 vssd1 vccd1 vccd1 _15566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 _15572_/Q vssd1 vssd1 vccd1 vccd1 hold2286/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08869_ _12380_/B _12445_/B vssd1 vssd1 vccd1 vccd1 _08912_/S sky130_fd_sc_hd__or2_2
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1552 hold1552/A vssd1 vssd1 vccd1 vccd1 input42/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2297 _15860_/Q vssd1 vssd1 vccd1 vccd1 hold2297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1563 _15618_/Q vssd1 vssd1 vccd1 vccd1 hold1563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 _15160_/X vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ hold5276/X _11198_/B _10899_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10900_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1585 _15561_/Q vssd1 vssd1 vccd1 vccd1 hold1585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1596 _08481_/X vssd1 vssd1 vccd1 vccd1 _15869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ _12267_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__or2_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10831_ hold3810/X _11095_/A2 _10830_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13550_ hold2020/X hold4321/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13551_/B sky130_fd_sc_hd__mux2_1
X_10762_ hold5591/X _11147_/B _10761_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ hold5/X _12509_/A2 _12507_/A3 _12500_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold6/A sky130_fd_sc_hd__o311a_1
XFILLER_0_165_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ hold2420/X _17614_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ hold5046/X _11168_/B _10692_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _10693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ hold887/X _15219_/B _15219_/Y _15030_/A vssd1 vssd1 vccd1 vccd1 hold888/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _12436_/A hold285/X vssd1 vssd1 vccd1 vccd1 _17309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _15205_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ hold3623/X _12267_/A _12362_/X vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14102_ _15229_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ hold4399/X _11801_/B _11313_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__o211a_1
X_15082_ hold3151/X _15113_/B _15081_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15082_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ hold4641/X _12288_/A _12293_/X vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_238_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ hold2834/X _14040_/B _14032_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14033_/X
+ sky130_fd_sc_hd__o211a_1
X_11245_ hold3948/X _11726_/B _11244_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11176_ _12340_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _16882_/D sky130_fd_sc_hd__nor2_1
XTAP_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10127_ hold3004/X hold4637/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _18300_/CLK _15984_/D vssd1 vssd1 vccd1 vccd1 hold712/A sky130_fd_sc_hd__dfxtp_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _17723_/CLK _17723_/D vssd1 vssd1 vccd1 vccd1 _17723_/Q sky130_fd_sc_hd__dfxtp_1
X_14935_ hold1695/X _14946_/B _14934_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _10058_/A _10070_/B _10190_/S vssd1 vssd1 vccd1 vccd1 _10058_/X sky130_fd_sc_hd__and3_1
XFILLER_0_234_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _17686_/CLK _17654_/D vssd1 vssd1 vccd1 vccd1 _17654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14866_ _15205_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_203_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16605_ _18225_/CLK _16605_/D vssd1 vssd1 vccd1 vccd1 _16605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13817_ _17726_/Q _13817_/B _13817_/C vssd1 vssd1 vccd1 vccd1 _13817_/X sky130_fd_sc_hd__and3_1
X_17585_ _17585_/CLK _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
X_14797_ hold3027/X _14828_/B _14796_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14797_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17299_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16536_ _17968_/CLK _16536_/D vssd1 vssd1 vccd1 vccd1 _16536_/Q sky130_fd_sc_hd__dfxtp_1
X_13748_ hold1992/X _17703_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16467_ _18378_/CLK _16467_/D vssd1 vssd1 vccd1 vccd1 _16467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13679_ hold2469/X hold4344/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18206_ _18232_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
X_15418_ hold235/X _09367_/A _15479_/B1 _17345_/Q vssd1 vssd1 vccd1 vccd1 _15418_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _18309_/CLK _16398_/D vssd1 vssd1 vccd1 vccd1 _16398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ _18233_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
X_15349_ hold899/X _09365_/B _09392_/C hold878/X _15348_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5807 hold5941/X vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5818 hold5944/X vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__buf_1
Xhold5829 hold5950/X vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold104 hold245/X vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18068_ _18068_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold148 hold7/X vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ hold4050/X _10004_/B _09909_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09910_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17019_ _17897_/CLK _17019_/D vssd1 vssd1 vccd1 vccd1 _17019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout606 _15488_/A2 vssd1 vssd1 vccd1 vccd1 _09392_/C sky130_fd_sc_hd__buf_6
X_09841_ hold3936/X _10007_/B _09840_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09841_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout617 _09354_/Y vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_238_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout628 _07824_/Y vssd1 vssd1 vccd1 vccd1 _15477_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_225_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout639 _12696_/A vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ hold5677/X _10070_/B _09771_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09772_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ hold292/X hold298/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__mux2_1
XFILLER_0_198_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08654_ _15324_/A hold548/X vssd1 vssd1 vccd1 vccd1 _15949_/D sky130_fd_sc_hd__and2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08585_ _15344_/A hold680/X vssd1 vssd1 vccd1 vccd1 _15916_/D sky130_fd_sc_hd__and2_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _15535_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ hold1057/X _09177_/A2 _09136_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _09137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_446_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09068_ _15509_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08019_ _15533_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__or2_1
Xhold660 hold660/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 hold671/A vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11030_ hold2919/X hold4553/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11031_/B sky130_fd_sc_hd__mux2_1
Xhold682 hold745/X vssd1 vssd1 vccd1 vccd1 hold746/A sky130_fd_sc_hd__buf_6
Xhold693 hold693/A vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2050 _09077_/X vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2061 _18434_/Q vssd1 vssd1 vccd1 vccd1 hold2061/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _15669_/Q vssd1 vssd1 vccd1 vccd1 hold2072/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2083 _15886_/Q vssd1 vssd1 vccd1 vccd1 hold2083/X sky130_fd_sc_hd__dlygate4sd3_1
X_12981_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _17503_/D sky130_fd_sc_hd__and2_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2094 _17998_/Q vssd1 vssd1 vccd1 vccd1 hold2094/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_232_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _14059_/X vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ _14774_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__nand2_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1371 _15634_/Q vssd1 vssd1 vccd1 vccd1 hold1371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1382 _09403_/X vssd1 vssd1 vccd1 vccd1 _16287_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ hold5419/X _12031_/A2 _11931_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11932_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _17995_/Q vssd1 vssd1 vccd1 vccd1 hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ hold2498/X _14666_/B _14650_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14651_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ hold4409/X _12365_/B _11862_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11863_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ hold1458/X _16762_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__mux2_1
X_13602_ _13734_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__or2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17370_ _17370_/CLK _17370_/D vssd1 vssd1 vccd1 vccd1 _17370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _15191_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__or2_1
X_11794_ _12367_/A _11794_/B vssd1 vssd1 vccd1 vccd1 _17088_/D sky130_fd_sc_hd__nor2_1
X_16321_ _16322_/CLK _16321_/D vssd1 vssd1 vccd1 vccd1 hold850/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10745_ hold1503/X hold4992/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__mux2_1
X_13533_ _13734_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _13533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ _13746_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__or2_1
X_16252_ _17431_/CLK _16252_/D vssd1 vssd1 vccd1 vccd1 _16252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10676_ hold1442/X hold4911/X _11159_/C vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15203_ _15203_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ hold379/X hold492/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ _13779_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__or2_1
X_16183_ _17479_/CLK _16183_/D vssd1 vssd1 vccd1 vccd1 _16183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ hold5996/X _15165_/B hold747/X _15066_/A vssd1 vssd1 vccd1 vccd1 hold748/A
+ sky130_fd_sc_hd__o211a_1
X_12346_ _13873_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _17272_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_187_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_116_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15065_ _15227_/A hold2479/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15066_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12277_ hold4475/X _13877_/B _12276_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12277_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _15523_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14016_/X sky130_fd_sc_hd__or2_1
X_11228_ _18424_/Q _16900_/Q _11711_/S vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ _16877_/Q _11159_/B _11159_/C vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__and3_1
XTAP_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _17286_/CLK _15967_/D vssd1 vssd1 vccd1 vccd1 hold537/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17706_ _17738_/CLK _17706_/D vssd1 vssd1 vccd1 vccd1 _17706_/Q sky130_fd_sc_hd__dfxtp_1
X_14918_ _14972_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14918_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15898_ _17344_/CLK _15898_/D vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__dfxtp_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17637_ _17701_/CLK _17637_/D vssd1 vssd1 vccd1 vccd1 _17637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14849_ hold874/X _14882_/B _14848_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 hold875/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08370_ _15539_/A hold2537/X hold134/X vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__mux2_1
X_17568_ _17696_/CLK _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ _18296_/CLK _16519_/D vssd1 vssd1 vccd1 vccd1 _16519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _17499_/CLK _17499_/D vssd1 vssd1 vccd1 vccd1 _17499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5604 _11410_/X vssd1 vssd1 vccd1 vccd1 _16960_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5615 _16802_/Q vssd1 vssd1 vccd1 vccd1 hold5615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5626 _10915_/X vssd1 vssd1 vccd1 vccd1 _16795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5637 _16983_/Q vssd1 vssd1 vccd1 vccd1 hold5637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4903 _16715_/Q vssd1 vssd1 vccd1 vccd1 hold4903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5648 _17047_/Q vssd1 vssd1 vccd1 vccd1 hold5648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5659 _17567_/Q vssd1 vssd1 vccd1 vccd1 hold5659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4914 _12103_/X vssd1 vssd1 vccd1 vccd1 _17191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4925 _16593_/Q vssd1 vssd1 vccd1 vccd1 hold4925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4936 _16559_/Q vssd1 vssd1 vccd1 vccd1 hold4936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4947 _12190_/X vssd1 vssd1 vccd1 vccd1 _17220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4958 _16565_/Q vssd1 vssd1 vccd1 vccd1 hold4958/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4969 _10393_/X vssd1 vssd1 vccd1 vccd1 _16621_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout403 _14338_/B vssd1 vssd1 vccd1 vccd1 _14336_/B sky130_fd_sc_hd__buf_8
Xfanout414 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14142_/B sky130_fd_sc_hd__buf_6
Xfanout425 hold123/X vssd1 vssd1 vccd1 vccd1 _13942_/S sky130_fd_sc_hd__clkbuf_8
Xfanout436 _13622_/S vssd1 vssd1 vccd1 vccd1 _12302_/C sky130_fd_sc_hd__buf_4
X_09824_ hold1232/X _16432_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__mux2_1
Xfanout447 _11150_/C vssd1 vssd1 vccd1 vccd1 _11711_/S sky130_fd_sc_hd__buf_4
XFILLER_0_226_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout458 _13847_/C vssd1 vssd1 vccd1 vccd1 _13871_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout469 _10025_/C vssd1 vssd1 vccd1 vccd1 _12368_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09755_ hold1787/X _16409_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09756_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_216_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08706_ _12408_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ hold2871/X hold5162/X _10190_/S vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08637_ hold402/X hold539/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__mux2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ hold568/X hold651/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__mux2_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08499_ hold1289/X _08486_/B _08498_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ _10533_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _11100_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ hold1159/X hold4927/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_280_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18214_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13180_ hold4664/X _13179_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_241_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ _10488_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12131_ hold1369/X hold3464/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12062_ hold1221/X hold3456/X _13868_/C vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__mux2_1
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11013_ _11115_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11013_/X sky130_fd_sc_hd__or2_1
X_16870_ _18039_/CLK _16870_/D vssd1 vssd1 vccd1 vccd1 _16870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _17732_/CLK _15821_/D vssd1 vssd1 vccd1 vccd1 hold663/A sky130_fd_sc_hd__dfxtp_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _17703_/CLK _15752_/D vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ hold1775/X hold3171/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__mux2_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 _15750_/Q vssd1 vssd1 vccd1 vccd1 hold1190/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ hold3116/X _14714_/B _14702_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14703_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ hold2072/X _17129_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15683_ _17775_/CLK _15683_/D vssd1 vssd1 vccd1 vccd1 _15683_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12895_ hold2395/X _17476_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__mux2_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17422_ _17422_/CLK _17422_/D vssd1 vssd1 vccd1 vccd1 _17422_/Q sky130_fd_sc_hd__dfxtp_1
X_14634_ _15189_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14634_/X sky130_fd_sc_hd__or2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11846_ hold1316/X hold3645/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11847_/B sky130_fd_sc_hd__mux2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17353_ _17515_/CLK _17353_/D vssd1 vssd1 vccd1 vccd1 _17353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _15189_/A _14557_/Y hold2088/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _14565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11777_ _17083_/Q _12317_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _11777_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _18405_/CLK hold896/X vssd1 vssd1 vccd1 vccd1 _16304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13516_ hold4247/X _13802_/B _13515_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10728_ _11124_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
X_17284_ _17284_/CLK _17284_/D vssd1 vssd1 vccd1 vccd1 hold704/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_368_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17734_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14496_ hold2814/X _14487_/B _14495_/X _12981_/A vssd1 vssd1 vccd1 vccd1 _14496_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16235_ _17429_/CLK _16235_/D vssd1 vssd1 vccd1 vccd1 _16235_/Q sky130_fd_sc_hd__dfxtp_1
X_13447_ hold5721/X _13829_/B _13446_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _11637_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13378_ hold3484/X _13847_/B _13377_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__o211a_1
X_16166_ _17879_/CLK _16166_/D vssd1 vssd1 vccd1 vccd1 _16166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15117_ hold559/X hold734/X vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__or2_1
X_12329_ _17267_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__and3_1
XFILLER_0_80_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16097_ _16097_/CLK _16097_/D vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3509 _17703_/Q vssd1 vssd1 vccd1 vccd1 hold3509/X sky130_fd_sc_hd__dlygate4sd3_1
X_15048_ _15052_/A _15048_/B vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__and2_1
XFILLER_0_177_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2808 _16224_/Q vssd1 vssd1 vccd1 vccd1 hold2808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2819 _18446_/Q vssd1 vssd1 vccd1 vccd1 hold2819/X sky130_fd_sc_hd__dlygate4sd3_1
X_07870_ hold2607/X _07869_/B _07869_/Y _08147_/A vssd1 vssd1 vccd1 vccd1 _07870_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16999_ _17877_/CLK _16999_/D vssd1 vssd1 vccd1 vccd1 _16999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09540_ _09918_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_84_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17161_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09471_ _09472_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__or2_1
Xclkbuf_6_41_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_41_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ hold1652/X _08433_/B _08421_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _08422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08353_ _08353_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08284_ hold202/X hold733/X vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__or2_4
XFILLER_0_73_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5401 _17261_/Q vssd1 vssd1 vccd1 vccd1 hold5401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5412 _11257_/X vssd1 vssd1 vccd1 vccd1 _16909_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5423 _17040_/Q vssd1 vssd1 vccd1 vccd1 hold5423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5434 _10141_/X vssd1 vssd1 vccd1 vccd1 _16537_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4700 _11163_/Y vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5445 _17275_/Q vssd1 vssd1 vccd1 vccd1 hold5445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4711 _16330_/Q vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5456 _12163_/X vssd1 vssd1 vccd1 vccd1 _17211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4722 _10486_/X vssd1 vssd1 vccd1 vccd1 _16652_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5467 _16797_/Q vssd1 vssd1 vccd1 vccd1 hold5467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4733 _16483_/Q vssd1 vssd1 vccd1 vccd1 hold4733/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5478 _10750_/X vssd1 vssd1 vccd1 vccd1 _16740_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4744 _09646_/X vssd1 vssd1 vccd1 vccd1 _16372_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5489 _17265_/Q vssd1 vssd1 vccd1 vccd1 hold5489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4755 _16373_/Q vssd1 vssd1 vccd1 vccd1 hold4755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4766 _09778_/X vssd1 vssd1 vccd1 vccd1 _16416_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout200 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__clkbuf_4
Xhold4777 _16513_/Q vssd1 vssd1 vccd1 vccd1 hold4777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout211 _09832_/A2 vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__buf_4
Xhold4788 _12312_/Y vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout222 _11192_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__buf_4
Xfanout233 _10565_/B vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__buf_4
Xhold4799 _16584_/Q vssd1 vssd1 vccd1 vccd1 hold4799/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout244 _10037_/B vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout255 _12024_/A vssd1 vssd1 vccd1 vccd1 _13794_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout266 _11139_/A vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__buf_2
XFILLER_0_236_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09807_ _11064_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__or2_1
Xfanout277 _13779_/A vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__buf_4
Xfanout288 _11679_/A vssd1 vssd1 vccd1 vccd1 _12057_/A sky130_fd_sc_hd__buf_4
Xfanout299 _09843_/A vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__buf_4
X_07999_ _14794_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _07999_/X sky130_fd_sc_hd__or2_1
XFILLER_0_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ _09984_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09669_ _10191_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__or2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _12246_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ hold3801/X _12679_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__mux2_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__or2_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ _14350_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _17972_/D sky130_fd_sc_hd__and2_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11562_ _11658_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_461_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10513_ hold4932/X _10631_/B _10512_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10513_/X
+ sky130_fd_sc_hd__o211a_1
X_13301_ _13300_/X hold3607/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14281_ hold2387/X _14266_/B _14280_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ _12219_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13232_ _13225_/X _13231_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__o21a_1
X_16020_ _17315_/CLK _16020_/D vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__dfxtp_1
X_10444_ hold5026/X _11180_/B _10443_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13163_ _13162_/X hold3583/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ hold5092/X _10571_/B _10374_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12114_ _12213_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13094_ _13094_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__or2_1
Xhold5990 _18016_/Q vssd1 vssd1 vccd1 vccd1 hold5990/X sky130_fd_sc_hd__dlygate4sd3_1
X_17971_ _17971_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12045_ _13773_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__or2_1
X_16922_ _17896_/CLK _16922_/D vssd1 vssd1 vccd1 vccd1 _16922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16853_ _18054_/CLK _16853_/D vssd1 vssd1 vccd1 vccd1 _16853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15804_ _17737_/CLK _15804_/D vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16784_ _17985_/CLK _16784_/D vssd1 vssd1 vccd1 vccd1 _16784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _14443_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13996_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15735_ _17738_/CLK _15735_/D vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12947_ hold3270/X _12946_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__mux2_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18455_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666_ _17200_/CLK _15666_/D vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ hold3299/X _12877_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17405_ _18455_/CLK _17405_/D vssd1 vssd1 vccd1 vccd1 _17405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ hold1676/X _14612_/B _14616_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14617_/X
+ sky130_fd_sc_hd__o211a_1
X_18385_ _18391_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _12213_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15597_ _17245_/CLK _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17344_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 _17336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14548_ hold2693/X _14541_/B _14547_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_131_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17267_ _17899_/CLK _17267_/D vssd1 vssd1 vccd1 vccd1 _17267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14479_ _15105_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16218_ _17878_/CLK _16218_/D vssd1 vssd1 vccd1 vccd1 _16218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _17198_/CLK _17198_/D vssd1 vssd1 vccd1 vccd1 _17198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4007 _09727_/X vssd1 vssd1 vccd1 vccd1 _16399_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16149_ _17508_/CLK _16149_/D vssd1 vssd1 vccd1 vccd1 _16149_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4018 _16785_/Q vssd1 vssd1 vccd1 vccd1 hold4018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4029 _10369_/X vssd1 vssd1 vccd1 vccd1 _16613_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3306 _17576_/Q vssd1 vssd1 vccd1 vccd1 hold3306/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3317 _17439_/Q vssd1 vssd1 vccd1 vccd1 hold3317/X sky130_fd_sc_hd__dlygate4sd3_1
X_08971_ hold568/X hold685/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3328 _17575_/Q vssd1 vssd1 vccd1 vccd1 hold3328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3339 _12776_/X vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2605 _15597_/Q vssd1 vssd1 vccd1 vccd1 hold2605/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2616 _15667_/Q vssd1 vssd1 vccd1 vccd1 hold2616/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _15545_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__nand2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2627 _09163_/X vssd1 vssd1 vccd1 vccd1 _16194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 _15736_/Q vssd1 vssd1 vccd1 vccd1 hold2638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 _08026_/X vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _17934_/Q vssd1 vssd1 vccd1 vccd1 hold1904/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1915 _14875_/X vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _14758_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__or2_1
Xhold1926 _14039_/X vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1937 _18197_/Q vssd1 vssd1 vccd1 vccd1 hold1937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1948 _15560_/X vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 _14289_/X vssd1 vssd1 vccd1 vccd1 _17942_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _18459_/Q vssd1 vssd1 vccd1 vccd1 _14556_/A sky130_fd_sc_hd__inv_2
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ hold3422/X _10025_/B _09522_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _09523_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ _09455_/B _09484_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _16311_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08405_ _15519_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_219_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18141_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09385_ hold5864/A _09342_/B _09342_/Y _09384_/X _12412_/A vssd1 vssd1 vccd1 vccd1
+ _09385_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_136_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08336_ hold1755/X _08336_/A2 _08335_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ hold2597/X _08268_/B _08266_/Y _13720_/C1 vssd1 vssd1 vccd1 vccd1 _08267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08198_ hold2436/X _08213_/B _08197_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5220 _17070_/Q vssd1 vssd1 vccd1 vccd1 hold5220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5231 _11590_/X vssd1 vssd1 vccd1 vccd1 _17020_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5242 _17071_/Q vssd1 vssd1 vccd1 vccd1 hold5242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5253 _09904_/X vssd1 vssd1 vccd1 vccd1 _16458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5264 _16813_/Q vssd1 vssd1 vccd1 vccd1 hold5264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5275 _12100_/X vssd1 vssd1 vccd1 vccd1 _17190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4530 _12247_/X vssd1 vssd1 vccd1 vccd1 _17239_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ hold1676/X hold3571/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__mux2_1
Xhold5286 _16867_/Q vssd1 vssd1 vccd1 vccd1 hold5286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4541 _17732_/Q vssd1 vssd1 vccd1 vccd1 hold4541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5297 _12220_/X vssd1 vssd1 vccd1 vccd1 _17230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4552 _12058_/X vssd1 vssd1 vccd1 vccd1 _17176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4563 _17700_/Q vssd1 vssd1 vccd1 vccd1 hold4563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4574 _15472_/X vssd1 vssd1 vccd1 vccd1 _15473_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4585 hold5817/X vssd1 vssd1 vccd1 vccd1 hold4585/X sky130_fd_sc_hd__buf_4
Xhold3840 _10138_/X vssd1 vssd1 vccd1 vccd1 _16536_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4596 _10038_/Y vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10091_ hold2109/X _16521_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__mux2_1
Xhold3851 _11220_/Y vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3862 _16931_/Q vssd1 vssd1 vccd1 vccd1 hold3862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3873 _10426_/X vssd1 vssd1 vccd1 vccd1 _16632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3884 _16842_/Q vssd1 vssd1 vccd1 vccd1 hold3884/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3895 _10768_/X vssd1 vssd1 vccd1 vccd1 _16746_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _17737_/Q _13880_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__and3_1
XFILLER_0_236_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12801_ _12810_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _17443_/D sky130_fd_sc_hd__and2_1
XFILLER_0_202_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10993_ hold4095/X _11095_/A2 _10992_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _10993_/X
+ sky130_fd_sc_hd__o211a_1
X_13781_ hold2555/X hold3490/X _13877_/C vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ hold1100/X _15507_/Y _15519_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _15520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12738_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _17420_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ hold654/X _15451_/A2 _09386_/D hold342/X _15446_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/D sky130_fd_sc_hd__a221o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12663_ _12738_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _17397_/D sky130_fd_sc_hd__and2_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ hold3118/X _14446_/A2 _14401_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14402_/X
+ sky130_fd_sc_hd__o211a_1
X_18170_ _18170_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_11614_ hold5036/X _12317_/B _11613_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11614_/X
+ sky130_fd_sc_hd__o211a_1
X_15382_ _15480_/A _15382_/B _15382_/C _15382_/D vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12594_ _12600_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _17374_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17121_ _17585_/CLK _17121_/D vssd1 vssd1 vccd1 vccd1 _17121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ hold2709/X hold756/X _14332_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ hold5334/X _11732_/B _11544_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _11545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17052_ _17265_/CLK _17052_/D vssd1 vssd1 vccd1 vccd1 _17052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14264_ _15105_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ hold5437/X _11762_/B _11475_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11476_/X
+ sky130_fd_sc_hd__o211a_1
X_16003_ _18408_/CLK _16003_/D vssd1 vssd1 vccd1 vccd1 hold775/A sky130_fd_sc_hd__dfxtp_1
X_10427_ hold1161/X _16633_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__mux2_1
X_13215_ _13311_/A1 _13213_/X _13214_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13215_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14195_ hold2737/X _14198_/B _14194_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ hold3143/X _16610_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _17569_/Q _17103_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13077_ _13076_/X hold4329/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__mux2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _18018_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
X_10289_ hold3006/X _16587_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12028_ hold5375/X _13862_/B _12027_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12028_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16905_ _17815_/CLK _16905_/D vssd1 vssd1 vccd1 vccd1 _16905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17885_ _17885_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16836_ _18071_/CLK _16836_/D vssd1 vssd1 vccd1 vccd1 _16836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _17968_/CLK _16767_/D vssd1 vssd1 vccd1 vccd1 _16767_/Q sky130_fd_sc_hd__dfxtp_1
X_13979_ hold2925/X _13986_/B _13978_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _13979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ _17253_/CLK _15718_/D vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_383_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17198_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16698_ _18222_/CLK _16698_/D vssd1 vssd1 vccd1 vccd1 _16698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18437_ _18453_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_312_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17971_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15649_ _17161_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09170_ _15553_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__or2_1
X_18368_ _18373_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ _13933_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__and2_1
X_17319_ _17320_/CLK hold114/X vssd1 vssd1 vccd1 vccd1 _17319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18299_ _18363_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08052_ hold999/X _08094_/B vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3103 _07957_/X vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3114 _18171_/Q vssd1 vssd1 vccd1 vccd1 hold3114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3125 _14414_/X vssd1 vssd1 vccd1 vccd1 _18003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3136 _17505_/Q vssd1 vssd1 vccd1 vccd1 hold3136/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3147 _18245_/Q vssd1 vssd1 vccd1 vccd1 hold3147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2402 _09213_/X vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08954_ _09053_/A hold191/X vssd1 vssd1 vccd1 vccd1 _16094_/D sky130_fd_sc_hd__and2_1
Xhold3158 _12530_/X vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2413 _17988_/Q vssd1 vssd1 vccd1 vccd1 hold2413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3169 _14933_/X vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _15681_/Q vssd1 vssd1 vccd1 vccd1 hold2424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 _14089_/X vssd1 vssd1 vccd1 vccd1 _17847_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1701 _17992_/Q vssd1 vssd1 vccd1 vccd1 hold1701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2446 _08237_/X vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07905_ hold2343/X _07924_/B _07904_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07905_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2457 _16273_/Q vssd1 vssd1 vccd1 vccd1 hold2457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1712 _17791_/Q vssd1 vssd1 vccd1 vccd1 hold1712/X sky130_fd_sc_hd__dlygate4sd3_1
X_08885_ _15344_/A hold890/X vssd1 vssd1 vccd1 vccd1 _16060_/D sky130_fd_sc_hd__and2_1
Xhold1723 hold1891/X vssd1 vssd1 vccd1 vccd1 hold1723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 _14075_/X vssd1 vssd1 vccd1 vccd1 _17840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _15144_/X vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2479 _18316_/Q vssd1 vssd1 vccd1 vccd1 hold2479/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1745 _08501_/X vssd1 vssd1 vccd1 vccd1 _15879_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 _08336_/X vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07836_ hold2880/X _07865_/B _07835_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _07836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1767 _15639_/Q vssd1 vssd1 vccd1 vccd1 hold1767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1778 _09423_/X vssd1 vssd1 vccd1 vccd1 _16297_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1789 _18106_/Q vssd1 vssd1 vccd1 vccd1 hold1789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09506_ hold1805/X _13078_/A _10004_/C vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _07785_/Y hold895/X _12412_/A _09436_/X vssd1 vssd1 vccd1 vccd1 hold896/A
+ sky130_fd_sc_hd__o211a_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09368_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08319_ _15543_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08319_/Y sky130_fd_sc_hd__nand2_1
X_09299_ _14910_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_60 hold746/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_71 _15203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 hold181/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ hold1119/X _16934_/Q _11711_/S vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__mux2_1
XANTENNA_93 hold746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11261_ hold2065/X hold4681/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5050 _16815_/Q vssd1 vssd1 vccd1 vccd1 hold5050/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5061 _10231_/X vssd1 vssd1 vccd1 vccd1 _16567_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10212_ _10524_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__or2_1
X_13000_ hold1919/X _07826_/A _13000_/S vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11192_ _11192_/A _11192_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__and3_1
Xhold5072 _17131_/Q vssd1 vssd1 vccd1 vccd1 hold5072/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5083 _10234_/X vssd1 vssd1 vccd1 vccd1 _16568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5094 _16482_/Q vssd1 vssd1 vccd1 vccd1 hold5094/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4360 _17048_/Q vssd1 vssd1 vccd1 vccd1 hold4360/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10143_ _10527_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4371 _12178_/X vssd1 vssd1 vccd1 vccd1 _17216_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4382 _17187_/Q vssd1 vssd1 vccd1 vccd1 hold4382/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4393 _17704_/Q vssd1 vssd1 vccd1 vccd1 hold4393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3670 _16929_/Q vssd1 vssd1 vccd1 vccd1 hold3670/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ hold1981/X _14952_/B _14950_/Y _15162_/C1 vssd1 vssd1 vccd1 vccd1 _14951_/X
+ sky130_fd_sc_hd__o211a_1
X_10074_ _13310_/A _10488_/A _10073_/X vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3681 _16481_/Q vssd1 vssd1 vccd1 vccd1 hold3681/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3692 _11175_/Y vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _14403_/A hold2065/X hold124/X vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__mux2_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2980 _15104_/X vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17670_ _17702_/CLK _17670_/D vssd1 vssd1 vccd1 vccd1 _17670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ _15221_/A _14882_/B vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__nand2_1
Xhold2991 _16161_/Q vssd1 vssd1 vccd1 vccd1 hold2991/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16621_ _18209_/CLK _16621_/D vssd1 vssd1 vccd1 vccd1 _16621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ hold5667/X _13698_/A _13832_/X vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16552_ _18108_/CLK _16552_/D vssd1 vssd1 vccd1 vccd1 _16552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ _13788_/A _13764_/B vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__or2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ hold2874/X hold5409/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15503_ hold525/X _18429_/Q hold691/X vssd1 vssd1 vccd1 vccd1 hold692/A sky130_fd_sc_hd__mux2_1
X_12715_ hold3035/X _17416_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16483_ _18266_/CLK _16483_/D vssd1 vssd1 vccd1 vccd1 _16483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _13779_/A _13695_/B vssd1 vssd1 vccd1 vccd1 _13695_/X sky130_fd_sc_hd__or2_1
XFILLER_0_210_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18222_ _18222_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15434_ _15482_/A _15434_/B vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ hold2566/X hold3468/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18153_ _18153_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ hold484/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ hold3045/X hold3159/X _12967_/S vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _17718_/CLK _17104_/D vssd1 vssd1 vccd1 vccd1 _17104_/Q sky130_fd_sc_hd__dfxtp_1
X_14316_ _15103_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__or2_1
X_18084_ _18208_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11528_ hold2725/X hold5062/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__mux2_1
X_15296_ _17333_/Q _15448_/B1 _15485_/B1 hold348/X vssd1 vssd1 vccd1 vccd1 _15296_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17035_ _18425_/CLK _17035_/D vssd1 vssd1 vccd1 vccd1 _17035_/Q sky130_fd_sc_hd__dfxtp_1
X_14247_ hold2317/X _14266_/B _14246_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14247_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11459_ hold1925/X hold4487/X _11594_/S vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_238_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14178_ _14517_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__or2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13129_ _13129_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__and2_1
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 hold1106/X vssd1 vssd1 vccd1 vccd1 hold1107/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_237_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17937_ _17960_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 hold1047/X vssd1 vssd1 vccd1 vccd1 hold1019/X sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _12424_/A hold770/X vssd1 vssd1 vccd1 vccd1 _15956_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17868_ _17900_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ _18052_/CLK _16819_/D vssd1 vssd1 vccd1 vccd1 _16819_/Q sky130_fd_sc_hd__dfxtp_1
X_17799_ _17860_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09222_ _15551_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ hold1614/X _09164_/B _09152_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _09153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08104_ _15509_/A hold1172/X hold240/X vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__mux2_1
X_09084_ _14984_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08035_ _15549_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08035_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 hold820/A vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold831 hold831/A vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold864 hold864/A vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 hold886/A vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 hold897/A vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ hold2947/X _16486_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2210 _15685_/Q vssd1 vssd1 vccd1 vccd1 hold2210/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2221 _16187_/Q vssd1 vssd1 vccd1 vccd1 hold2221/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2232 _08491_/X vssd1 vssd1 vccd1 vccd1 _15874_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08937_ hold312/X hold549/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold550/A sky130_fd_sc_hd__mux2_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2243 _09203_/X vssd1 vssd1 vccd1 vccd1 _16213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_0_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2254 _16196_/Q vssd1 vssd1 vccd1 vccd1 hold2254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1520 _14887_/X vssd1 vssd1 vccd1 vccd1 _18230_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2265 _17933_/Q vssd1 vssd1 vccd1 vccd1 hold2265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2276 _17828_/Q vssd1 vssd1 vccd1 vccd1 hold2276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 _17763_/Q vssd1 vssd1 vccd1 vccd1 hold1531/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1542 _15644_/Q vssd1 vssd1 vccd1 vccd1 hold1542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 _07854_/X vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ _17520_/Q _08868_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1553 input42/X vssd1 vssd1 vccd1 vccd1 hold1553/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2298 _08463_/X vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _07951_/X vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1575 _15868_/Q vssd1 vssd1 vccd1 vccd1 hold1575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_234_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18225_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07819_ _15559_/A _15231_/A vssd1 vssd1 vccd1 vccd1 _09495_/C sky130_fd_sc_hd__nand2_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1586 _07832_/X vssd1 vssd1 vccd1 vccd1 _15561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _15867_/Q vssd1 vssd1 vccd1 vccd1 hold1597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08799_ hold312/X hold584/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold585/A sky130_fd_sc_hd__mux2_1
XFILLER_0_197_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _10830_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10761_ _11052_/A _10761_/B vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _17343_/Q _12500_/B vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13480_ hold5282/X _13817_/B _13479_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13480_/X
+ sky130_fd_sc_hd__o211a_1
X_10692_ _11070_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__or2_1
X_12431_ hold222/X hold284/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ hold1571/X _15165_/B _15149_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15150_/X
+ sky130_fd_sc_hd__o211a_1
X_12362_ _17278_/Q _13871_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ hold2776/X _14107_/A2 _14100_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11706_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__or2_1
X_15081_ _15189_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ _17255_/Q _12293_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__and3_1
XFILLER_0_132_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14032_ _15105_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__or2_1
X_11244_ _11631_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11175_ hold3691/X _11115_/A _11174_/X vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4190 _11038_/X vssd1 vssd1 vccd1 vccd1 _16836_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10126_ hold4873/X _10625_/B _10125_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10126_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15983_ _16127_/CLK _15983_/D vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _17722_/CLK _17722_/D vssd1 vssd1 vccd1 vccd1 _17722_/Q sky130_fd_sc_hd__dfxtp_1
X_10057_ _10603_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _16509_/D sky130_fd_sc_hd__nor2_1
X_14934_ _15203_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__or2_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _17747_/CLK _17653_/D vssd1 vssd1 vccd1 vccd1 _17653_/Q sky130_fd_sc_hd__dfxtp_1
X_14865_ hold2967/X _14880_/B _14864_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14865_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _18222_/CLK _16604_/D vssd1 vssd1 vccd1 vccd1 _16604_/Q sky130_fd_sc_hd__dfxtp_1
X_13816_ _13825_/A _13816_/B vssd1 vssd1 vccd1 vccd1 _17725_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_230_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17584_ _17712_/CLK _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
X_14796_ _15189_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14796_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16535_ _18123_/CLK _16535_/D vssd1 vssd1 vccd1 vccd1 _16535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13747_ hold4287/X _13847_/B _13746_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _11139_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16466_ _18377_/CLK _16466_/D vssd1 vssd1 vccd1 vccd1 _16466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ hold3511/X _13777_/A2 _13677_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13678_/X
+ sky130_fd_sc_hd__o211a_1
X_18205_ _18205_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15417_ hold190/X _09392_/B _09392_/C hold306/X vssd1 vssd1 vccd1 vccd1 _15417_/X
+ sky130_fd_sc_hd__a22o_1
X_12629_ hold3341/X _12628_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16397_ _18396_/CLK _16397_/D vssd1 vssd1 vccd1 vccd1 _16397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18136_ _18214_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15348_ hold834/X _09386_/A _15451_/A2 hold868/X vssd1 vssd1 vccd1 vccd1 _15348_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5808 output91/X vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_12
Xhold5819 output93/X vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18067_ _18067_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 hold37/X vssd1 vssd1 vccd1 vccd1 input10/A sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ hold374/X _15485_/A2 _15488_/A2 hold449/X _15278_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold138 hold10/X vssd1 vssd1 vccd1 vccd1 input25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 input29/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__buf_1
X_17018_ _17896_/CLK _17018_/D vssd1 vssd1 vccd1 vccd1 _17018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _09936_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__or2_1
Xfanout607 _09363_/Y vssd1 vssd1 vccd1 vccd1 _15488_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_10_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 _09351_/Y vssd1 vssd1 vccd1 vccd1 _15486_/A2 sky130_fd_sc_hd__buf_6
Xfanout629 _07824_/Y vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09771_ _10191_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _12408_/A hold194/X vssd1 vssd1 vccd1 vccd1 _15982_/D sky130_fd_sc_hd__and2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08653_ hold145/X hold547/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold548/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ hold210/X hold679/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold680/A sky130_fd_sc_hd__mux2_1
XFILLER_0_77_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09205_ hold2665/X _09218_/B _09204_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _09205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ _15519_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09067_ _15182_/A hold533/A vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__or2_2
XFILLER_0_124_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08018_ hold2411/X _08029_/B _08017_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _08018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 hold650/A vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 hold661/A vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 hold672/A vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 hold683/A vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold694/A vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _10467_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_415_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_1376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2040 _18448_/Q vssd1 vssd1 vccd1 vccd1 hold2040/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 _15741_/Q vssd1 vssd1 vccd1 vccd1 hold2051/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2062 _15516_/X vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2073 _08059_/X vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12980_ hold3219/X _12979_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_239_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2084 _08518_/X vssd1 vssd1 vccd1 vccd1 _15886_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 _15568_/Q vssd1 vssd1 vccd1 vccd1 hold1350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2095 _14404_/X vssd1 vssd1 vccd1 vccd1 _17998_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _17829_/Q vssd1 vssd1 vccd1 vccd1 hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _12261_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__or2_1
Xhold1372 _07983_/X vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 hold6050/X vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__buf_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _14398_/X vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14758_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__or2_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _12246_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11862_/X sky130_fd_sc_hd__or2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ hold2070/X _17654_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10813_ hold5451/X _11210_/B _10812_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ hold3236/X _14612_/B _14580_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14581_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ hold3685/X _11706_/A _11792_/X vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ _16320_/CLK _16320_/D vssd1 vssd1 vccd1 vccd1 _16320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13532_ hold2379/X hold5697/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ hold5563/X _11768_/B _10743_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _10744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16251_ _18455_/CLK _16251_/D vssd1 vssd1 vccd1 vccd1 _16251_/Q sky130_fd_sc_hd__dfxtp_1
X_13463_ hold2128/X hold3529/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__mux2_1
X_10675_ hold5535/X _11156_/B _10674_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _10675_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ hold3207/X _15221_/B _15201_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ _12426_/A _12414_/B vssd1 vssd1 vccd1 vccd1 _17300_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16182_ _17507_/CLK _16182_/D vssd1 vssd1 vccd1 vccd1 _16182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13394_ hold2231/X hold3312/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15133_ hold746/X _15171_/B vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__or2_1
X_12345_ hold3825/X _12057_/A _12344_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ _15064_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__and2_1
XFILLER_0_239_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12276_ _13782_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ hold2306/X _14040_/B _14014_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11227_ _12367_/A _11227_/B vssd1 vssd1 vccd1 vccd1 _16899_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_120_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11158_ _11158_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _16876_/D sky130_fd_sc_hd__nor2_1
XTAP_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ hold2291/X hold3553/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__mux2_1
X_15966_ _17293_/CLK _15966_/D vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
X_11089_ _11183_/A _11095_/A2 _11088_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14917_ hold1591/X _14952_/B _14916_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14917_/X
+ sky130_fd_sc_hd__o211a_1
X_17705_ _17737_/CLK _17705_/D vssd1 vssd1 vccd1 vccd1 _17705_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _16148_/CLK _15897_/D vssd1 vssd1 vccd1 vccd1 hold618/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_31_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_31_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14848_ hold746/X _14894_/B vssd1 vssd1 vccd1 vccd1 _14848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17636_ _17700_/CLK _17636_/D vssd1 vssd1 vccd1 vccd1 _17636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17567_ _17677_/CLK _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
X_14779_ hold1859/X _14772_/B _14778_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14779_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ _18234_/CLK _16518_/D vssd1 vssd1 vccd1 vccd1 _16518_/Q sky130_fd_sc_hd__dfxtp_1
X_17498_ _17499_/CLK _17498_/D vssd1 vssd1 vccd1 vccd1 _17498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16449_ _18394_/CLK _16449_/D vssd1 vssd1 vccd1 vccd1 _16449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18119_ _18175_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5605 _17074_/Q vssd1 vssd1 vccd1 vccd1 hold5605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5616 _10840_/X vssd1 vssd1 vccd1 vccd1 _16770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5627 _17042_/Q vssd1 vssd1 vccd1 vccd1 hold5627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5638 _11383_/X vssd1 vssd1 vccd1 vccd1 _16951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4904 _11154_/Y vssd1 vssd1 vccd1 vccd1 _11155_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5649 _11575_/X vssd1 vssd1 vccd1 vccd1 _17015_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4915 _17192_/Q vssd1 vssd1 vccd1 vccd1 hold4915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4926 _10213_/X vssd1 vssd1 vccd1 vccd1 _16561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4937 _10111_/X vssd1 vssd1 vccd1 vccd1 _16527_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4948 _16338_/Q vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4959 _10129_/X vssd1 vssd1 vccd1 vccd1 _16533_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout404 hold755/X vssd1 vssd1 vccd1 vccd1 hold756/A sky130_fd_sc_hd__buf_6
XFILLER_0_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout415 _14104_/B vssd1 vssd1 vccd1 vccd1 _14106_/B sky130_fd_sc_hd__buf_8
Xfanout426 _13307_/S vssd1 vssd1 vccd1 vccd1 _13251_/S sky130_fd_sc_hd__clkbuf_16
X_09823_ hold3976/X _10010_/B _09822_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09823_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout437 _13817_/C vssd1 vssd1 vccd1 vccd1 _13829_/C sky130_fd_sc_hd__buf_6
XFILLER_0_225_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout448 _11150_/C vssd1 vssd1 vccd1 vccd1 _11726_/C sky130_fd_sc_hd__clkbuf_8
Xfanout459 _13847_/C vssd1 vssd1 vccd1 vccd1 _13841_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09754_ hold5038/X _11177_/B _09753_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ hold353/X hold418/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08706_/B sky130_fd_sc_hd__mux2_1
X_09685_ hold4783/X _10565_/B _09684_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09685_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _15364_/A _08636_/B vssd1 vssd1 vccd1 vccd1 _15940_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08567_ _15364_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _15907_/D sky130_fd_sc_hd__and2_1
XFILLER_0_232_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08498_ _14443_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ hold2115/X _16644_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09119_ hold1919/X _09119_/A2 _09118_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09119_/X
+ sky130_fd_sc_hd__o211a_1
X_10391_ hold2516/X _16621_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ hold5272/X _13798_/A2 _12129_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12061_ hold3446/X _13868_/B _12060_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold480 hold480/A vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11012_ hold3220/X _16828_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _11013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15820_ _17667_/CLK _15820_/D vssd1 vssd1 vccd1 vccd1 _15820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15751_ _17702_/CLK _15751_/D vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _12969_/A _12963_/B vssd1 vssd1 vccd1 vccd1 _17497_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _13008_/X vssd1 vssd1 vccd1 vccd1 _17512_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14988_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14702_/X sky130_fd_sc_hd__or2_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 _08231_/X vssd1 vssd1 vccd1 vccd1 _15750_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ hold4972/X _13811_/B _11913_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _17210_/CLK _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12894_ _12894_/A _12894_/B vssd1 vssd1 vccd1 vccd1 _17474_/D sky130_fd_sc_hd__and2_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17422_/CLK _17421_/D vssd1 vssd1 vccd1 vccd1 _17421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14633_ hold1855/X _14666_/B _14632_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14633_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11845_ hold5116/X _12314_/B _11844_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17352_ _17515_/CLK _17352_/D vssd1 vssd1 vccd1 vccd1 _17352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ hold690/X _14573_/B hold2087/X vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__a21o_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12367_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _17082_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_56_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16322_/CLK hold851/X vssd1 vssd1 vccd1 vccd1 _16303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ _13713_/A _13515_/B vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__or2_1
X_17283_ _17283_/CLK _17283_/D vssd1 vssd1 vccd1 vccd1 _17283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10727_ hold1904/X _16733_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__mux2_1
X_14495_ _15229_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14495_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16234_ _17429_/CLK _16234_/D vssd1 vssd1 vccd1 vccd1 _16234_/Q sky130_fd_sc_hd__dfxtp_1
X_13446_ _13734_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__or2_1
X_10658_ hold1895/X hold3438/X _11729_/C vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _17879_/CLK _16165_/D vssd1 vssd1 vccd1 vccd1 _16165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ _13776_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _13377_/X sky130_fd_sc_hd__or2_1
X_10589_ _16687_/Q _10649_/B _10589_/C vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ hold2308/X _15111_/B _15115_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15116_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12328_ _13873_/A _12328_/B vssd1 vssd1 vccd1 vccd1 _17266_/D sky130_fd_sc_hd__nor2_1
X_16096_ _17304_/CLK _16096_/D vssd1 vssd1 vccd1 vccd1 hold783/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_337_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17153_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _15535_/A hold1313/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15048_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_220_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12259_ hold5445/X _12353_/B _12258_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2809 _09225_/X vssd1 vssd1 vccd1 vccd1 _16224_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16998_ _17876_/CLK _16998_/D vssd1 vssd1 vccd1 vccd1 _16998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15949_ _18402_/CLK _15949_/D vssd1 vssd1 vccd1 vccd1 hold547/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09470_ _09471_/B _09484_/B _09470_/C vssd1 vssd1 vccd1 vccd1 _16317_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08421_ _14529_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17619_ _17683_/CLK _17619_/D vssd1 vssd1 vccd1 vccd1 _17619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08352_ _15521_/A hold2037/X hold134/X vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18017_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ hold203/X hold733/X vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5402 _12217_/X vssd1 vssd1 vccd1 vccd1 _17229_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5413 _17220_/Q vssd1 vssd1 vccd1 vccd1 hold5413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5424 _11554_/X vssd1 vssd1 vccd1 vccd1 _17008_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5435 _17211_/Q vssd1 vssd1 vccd1 vccd1 hold5435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4701 _16537_/Q vssd1 vssd1 vccd1 vccd1 hold4701/X sky130_fd_sc_hd__buf_1
Xhold5446 _12259_/X vssd1 vssd1 vccd1 vccd1 _17243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4712 _09999_/Y vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5457 _16985_/Q vssd1 vssd1 vccd1 vccd1 hold5457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4723 _16419_/Q vssd1 vssd1 vccd1 vccd1 hold4723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5468 _10825_/X vssd1 vssd1 vccd1 vccd1 _16765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4734 _09883_/X vssd1 vssd1 vccd1 vccd1 _16451_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5479 _16804_/Q vssd1 vssd1 vccd1 vccd1 hold5479/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4745 _16682_/Q vssd1 vssd1 vccd1 vccd1 hold4745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4756 _09553_/X vssd1 vssd1 vccd1 vccd1 _16341_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4767 _16413_/Q vssd1 vssd1 vccd1 vccd1 hold4767/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout201 _11584_/A2 vssd1 vssd1 vccd1 vccd1 _12344_/B sky130_fd_sc_hd__buf_4
Xhold4778 _09973_/X vssd1 vssd1 vccd1 vccd1 _16481_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout212 _09832_/A2 vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4789 _16574_/Q vssd1 vssd1 vccd1 vccd1 hold4789/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout223 _10468_/A2 vssd1 vssd1 vccd1 vccd1 _11192_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout234 _10565_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__buf_4
Xfanout245 fanout246/X vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__buf_4
Xfanout256 _12024_/A vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__buf_4
X_09806_ hold988/X _16426_/Q _11159_/C vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__mux2_1
Xfanout267 _11070_/A vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__buf_4
XFILLER_0_214_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout278 _13779_/A vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__buf_4
X_07998_ hold1485/X _08033_/B _07997_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07998_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout289 _11679_/A vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__buf_4
XFILLER_0_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09737_ hold2273/X hold3359/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ hold1318/X hold5661/X _10190_/S vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ hold98/X hold667/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__mux2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ hold1841/X _16357_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__mux2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11630_ hold2860/X _17034_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11561_ hold1759/X _17011_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ hold4919/X _13299_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _10536_/A _10512_/B vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ _14782_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ hold2713/X hold3904/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _13311_/A1 _13229_/X _13230_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13231_/X
+ sky130_fd_sc_hd__o211a_1
X_10443_ _10830_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13162_ _17571_/Q _17105_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__mux2_1
X_10374_ _10560_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_430_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17686_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ hold2504/X hold5010/X _12308_/C vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5980 _18344_/Q vssd1 vssd1 vccd1 vccd1 hold5980/X sky130_fd_sc_hd__dlygate4sd3_1
X_13093_ _13092_/X hold4634/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__mux2_1
Xhold5991 _15842_/Q vssd1 vssd1 vccd1 vccd1 hold5991/X sky130_fd_sc_hd__dlygate4sd3_1
X_17970_ _17970_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
X_12044_ hold1258/X hold4233/X _13868_/C vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__mux2_1
X_16921_ _17767_/CLK _16921_/D vssd1 vssd1 vccd1 vccd1 _16921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16852_ _18053_/CLK _16852_/D vssd1 vssd1 vccd1 vccd1 _16852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout790 _13935_/A vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_4
XFILLER_0_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _17650_/CLK _15803_/D vssd1 vssd1 vccd1 vccd1 _15803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16783_ _18016_/CLK _16783_/D vssd1 vssd1 vccd1 vccd1 _16783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13995_ hold2430/X _13995_/A2 _13994_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _13995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15734_ _17737_/CLK _15734_/D vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ hold1123/X hold3256/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _18453_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
X_15665_ _17253_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ hold2603/X hold3288/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _15225_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14616_/X sky130_fd_sc_hd__or2_1
X_17404_ _18453_/CLK _17404_/D vssd1 vssd1 vccd1 vccd1 _17404_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _18384_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11828_ hold1023/X hold4645/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15596_ _17244_/CLK _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17335_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 _17335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14726_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _17077_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__and3_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _17266_/CLK _17266_/D vssd1 vssd1 vccd1 vccd1 _17266_/Q sky130_fd_sc_hd__dfxtp_1
X_14478_ hold3036/X _14482_/A2 _14477_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14478_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16217_ _17257_/CLK _16217_/D vssd1 vssd1 vccd1 vccd1 _16217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ hold4044/X _13802_/B _13428_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17197_ _17244_/CLK _17197_/D vssd1 vssd1 vccd1 vccd1 _17197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _16148_/CLK _16148_/D vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__dfxtp_1
Xhold4008 _16704_/Q vssd1 vssd1 vccd1 vccd1 hold4008/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_171_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4019 _10789_/X vssd1 vssd1 vccd1 vccd1 _16753_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08970_ _15324_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _16102_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18406_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _18401_/CLK _16079_/D vssd1 vssd1 vccd1 vccd1 hold464/A sky130_fd_sc_hd__dfxtp_1
Xhold3307 _13848_/Y vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3318 _12788_/X vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3329 _13845_/Y vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2606 _07907_/X vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07921_ hold2021/X _07924_/B _07920_/Y _13905_/A vssd1 vssd1 vccd1 vccd1 _07921_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2617 _08055_/X vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 _18342_/Q vssd1 vssd1 vccd1 vccd1 hold2628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2639 _08200_/X vssd1 vssd1 vccd1 vccd1 _15736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 _14271_/X vssd1 vssd1 vccd1 vccd1 _17934_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07852_ hold2969/X _07865_/B _07851_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _07852_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1916 _17761_/Q vssd1 vssd1 vccd1 vccd1 hold1916/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1927 _18118_/Q vssd1 vssd1 vccd1 vccd1 hold1927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 _14819_/X vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1949 _18428_/Q vssd1 vssd1 vccd1 vccd1 hold1949/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 input1/A vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07783_ hold469/X vssd1 vssd1 vccd1 vccd1 _07783_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09522_ _09984_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09453_ _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09455_/B sky130_fd_sc_hd__and3_1
XFILLER_0_56_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ hold2098/X _08440_/A2 _08403_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08404_/X
+ sky130_fd_sc_hd__o211a_1
X_09384_ hold630/X _15483_/B _09383_/X _18458_/Q vssd1 vssd1 vccd1 vccd1 _09384_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08335_ _14894_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08266_ _15545_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_259_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18036_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08197_ _14758_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08197_/X sky130_fd_sc_hd__or2_1
Xhold5210 _16613_/Q vssd1 vssd1 vccd1 vccd1 hold5210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5221 _11644_/X vssd1 vssd1 vccd1 vccd1 _17038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5232 _17126_/Q vssd1 vssd1 vccd1 vccd1 hold5232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5243 _11647_/X vssd1 vssd1 vccd1 vccd1 _17039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5254 _17167_/Q vssd1 vssd1 vccd1 vccd1 hold5254/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5265 _10873_/X vssd1 vssd1 vccd1 vccd1 _16781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4520 _11887_/X vssd1 vssd1 vccd1 vccd1 _17119_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4531 _16865_/Q vssd1 vssd1 vccd1 vccd1 hold4531/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5276 _16822_/Q vssd1 vssd1 vccd1 vccd1 hold5276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5287 _11035_/X vssd1 vssd1 vccd1 vccd1 _16835_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4542 _13741_/X vssd1 vssd1 vccd1 vccd1 _17700_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4553 _16834_/Q vssd1 vssd1 vccd1 vccd1 hold4553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5298 _17591_/Q vssd1 vssd1 vccd1 vccd1 hold5298/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4564 _13645_/X vssd1 vssd1 vccd1 vccd1 _17668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4575 _17676_/Q vssd1 vssd1 vccd1 vccd1 hold4575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3830 _11230_/X vssd1 vssd1 vccd1 vccd1 _16900_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10090_ hold4901/X _10598_/B _10089_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _10090_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4586 _15313_/X vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3841 _16821_/Q vssd1 vssd1 vccd1 vccd1 hold3841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4597 _16341_/Q vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3852 _16930_/Q vssd1 vssd1 vccd1 vccd1 hold3852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3863 _11802_/Y vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3874 _16609_/Q vssd1 vssd1 vccd1 vccd1 hold3874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3885 _10960_/X vssd1 vssd1 vccd1 vccd1 _16810_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3896 _16002_/Q vssd1 vssd1 vccd1 vccd1 _15325_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ hold3302/X _12799_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12801_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_187_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ hold3500/X _13886_/B _13779_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13780_/X
+ sky130_fd_sc_hd__o211a_1
X_10992_ _11094_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ hold3197/X _12730_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12731_/X sky130_fd_sc_hd__mux2_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ hold793/X _09365_/B _15485_/B1 hold543/X _15448_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_128_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ hold3521/X _12661_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _15189_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14401_/X sky130_fd_sc_hd__or2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11613_ _12285_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__or2_1
X_15381_ _16302_/Q _09362_/A _09392_/B hold739/X _15380_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_182_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ hold3230/X _12592_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12593_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17120_ _17280_/CLK _17120_/D vssd1 vssd1 vccd1 vccd1 _17120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ _14726_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11544_ _11553_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17051_ _17897_/CLK _17051_/D vssd1 vssd1 vccd1 vccd1 _17051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14263_ hold3059/X _14272_/B _14262_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ _11667_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16002_ _18407_/CLK _16002_/D vssd1 vssd1 vccd1 vccd1 _16002_/Q sky130_fd_sc_hd__dfxtp_1
X_13214_ _13214_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13214_/X sky130_fd_sc_hd__or2_1
X_10426_ hold3872/X _11095_/A2 _10425_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ _15539_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14194_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ _13145_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10357_ hold3956/X _10646_/B _10356_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ hold3438/X _13075_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__mux2_2
X_17953_ _17985_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
X_10288_ hold4859/X _11177_/B _10287_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12027_ _12261_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__or2_1
X_16904_ _17814_/CLK _16904_/D vssd1 vssd1 vccd1 vccd1 _16904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17884_ _17884_/CLK _17884_/D vssd1 vssd1 vccd1 vccd1 _17884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ _18036_/CLK _16835_/D vssd1 vssd1 vccd1 vccd1 _16835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13978_ _15105_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__or2_1
X_16766_ _17999_/CLK _16766_/D vssd1 vssd1 vccd1 vccd1 _16766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15717_ _17164_/CLK _15717_/D vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfxtp_1
X_12929_ hold3264/X _12928_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__mux2_1
X_16697_ _18221_/CLK _16697_/D vssd1 vssd1 vccd1 vccd1 _16697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18436_ _18436_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
X_15648_ _17160_/CLK hold983/X vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18367_ _18367_/CLK hold503/X vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ _17775_/CLK _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08120_ _15525_/A hold2965/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__mux2_1
X_17318_ _17320_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 _17318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_352_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17748_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18298_ _18362_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08051_ hold1243/X _08097_/A2 _08050_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08051_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17249_ _17585_/CLK _17249_/D vssd1 vssd1 vccd1 vccd1 _17249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3104 _18060_/Q vssd1 vssd1 vccd1 vccd1 hold3104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3115 _14765_/X vssd1 vssd1 vccd1 vccd1 _18171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3126 _16339_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_110_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ hold163/X hold190/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__mux2_1
Xhold3137 _12986_/X vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3148 _14921_/X vssd1 vssd1 vccd1 vccd1 _18245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2403 _15629_/Q vssd1 vssd1 vccd1 vccd1 hold2403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3159 _17370_/Q vssd1 vssd1 vccd1 vccd1 hold3159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 _17816_/Q vssd1 vssd1 vccd1 vccd1 hold2414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _08083_/X vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2436 _15735_/Q vssd1 vssd1 vccd1 vccd1 hold2436/X sky130_fd_sc_hd__dlygate4sd3_1
X_07904_ _14862_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1702 _18266_/Q vssd1 vssd1 vccd1 vccd1 hold1702/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ hold596/X hold889/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold890/A sky130_fd_sc_hd__mux2_1
Xhold2447 _18098_/Q vssd1 vssd1 vccd1 vccd1 hold2447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 _09326_/X vssd1 vssd1 vccd1 vccd1 _16273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 _13973_/X vssd1 vssd1 vccd1 vccd1 _17791_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2469 _15761_/Q vssd1 vssd1 vccd1 vccd1 hold2469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 hold1724/A vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__buf_12
Xhold1735 _15872_/Q vssd1 vssd1 vccd1 vccd1 hold1735/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1746 _15612_/Q vssd1 vssd1 vccd1 vccd1 hold1746/X sky130_fd_sc_hd__dlygate4sd3_1
X_07835_ _15513_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07835_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1757 _18103_/Q vssd1 vssd1 vccd1 vccd1 hold1757/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1768 _07996_/X vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 _16267_/Q vssd1 vssd1 vccd1 vccd1 hold1779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ hold3452/X _10025_/B _09504_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _09505_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ hold819/X _16304_/Q vssd1 vssd1 vccd1 vccd1 _09436_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09367_ _09367_/A _09386_/D vssd1 vssd1 vccd1 vccd1 _09369_/D sky130_fd_sc_hd__or2_1
XFILLER_0_30_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08318_ hold2315/X _08323_/B _08317_/Y _12657_/A vssd1 vssd1 vccd1 vccd1 _08318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09298_ hold1325/X _09338_/A2 _09297_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09298_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_50 _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_61 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_83 hold181/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ hold2375/X _08263_/A2 _08248_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _08249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_94 _15173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ hold5200/X _11738_/B _11259_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5040 _16454_/Q vssd1 vssd1 vccd1 vccd1 hold5040/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10211_ hold3055/X _16561_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__mux2_1
Xhold5051 _10879_/X vssd1 vssd1 vccd1 vccd1 _16783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5062 _17000_/Q vssd1 vssd1 vccd1 vccd1 hold5062/X sky130_fd_sc_hd__dlygate4sd3_1
X_11191_ _11218_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _16887_/D sky130_fd_sc_hd__nor2_1
Xhold5073 _11827_/X vssd1 vssd1 vccd1 vccd1 _17099_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5084 _16881_/Q vssd1 vssd1 vccd1 vccd1 hold5084/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4350 _17049_/Q vssd1 vssd1 vccd1 vccd1 hold4350/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5095 _09880_/X vssd1 vssd1 vccd1 vccd1 _16450_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10142_ hold2955/X hold3555/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__mux2_1
Xhold4361 _11578_/X vssd1 vssd1 vccd1 vccd1 _17016_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4372 _17683_/Q vssd1 vssd1 vccd1 vccd1 hold4372/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4383 _11995_/X vssd1 vssd1 vccd1 vccd1 _17155_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4394 _13657_/X vssd1 vssd1 vccd1 vccd1 _17672_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3660 _10093_/X vssd1 vssd1 vccd1 vccd1 _16521_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _15004_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14950_/Y sky130_fd_sc_hd__nand2_1
X_10073_ _16515_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__and3_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3671 _11796_/Y vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3682 _09877_/X vssd1 vssd1 vccd1 vccd1 _16449_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3693 _17416_/Q vssd1 vssd1 vccd1 vccd1 hold3693/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2970 _07852_/X vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13901_ _14378_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _17756_/D sky130_fd_sc_hd__and2_1
X_14881_ hold1970/X _14880_/B _14880_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2981 _18267_/Q vssd1 vssd1 vccd1 vccd1 hold2981/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2992 _09093_/X vssd1 vssd1 vccd1 vccd1 _16161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16620_ _18176_/CLK _16620_/D vssd1 vssd1 vccd1 vccd1 _16620_/Q sky130_fd_sc_hd__dfxtp_1
X_13832_ _17731_/Q _13832_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__and3_1
XFILLER_0_199_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16551_ _18263_/CLK _16551_/D vssd1 vssd1 vccd1 vccd1 _16551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ hold1628/X _17708_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10975_ hold3804/X _11168_/B _10974_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _10975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12714_ _12759_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _17414_/D sky130_fd_sc_hd__and2_1
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__and2_1
XFILLER_0_214_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ _18265_/CLK _16482_/D vssd1 vssd1 vccd1 vccd1 _16482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ hold2391/X hold3519/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18221_ _18221_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_15433_ _15481_/A1 _15425_/X _15432_/X _15481_/B1 _18417_/Q vssd1 vssd1 vccd1 vccd1
+ _15433_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_194_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ _12654_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _17391_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18152_ _18152_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_15364_ _15364_/A _15364_/B vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12576_ _12969_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _17368_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17103_ _17769_/CLK _17103_/D vssd1 vssd1 vccd1 vccd1 _17103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14315_ hold1511/X hold756/X _14314_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14315_/X
+ sky130_fd_sc_hd__o211a_1
X_18083_ _18223_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
X_11527_ hold5228/X _12299_/B _11526_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11527_/X
+ sky130_fd_sc_hd__o211a_1
X_15295_ hold842/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17034_ _17879_/CLK _17034_/D vssd1 vssd1 vccd1 vccd1 _17034_/Q sky130_fd_sc_hd__dfxtp_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ _14246_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ hold5246/X _11732_/B _11457_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10409_ hold1908/X hold3972/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14177_ hold2329/X _14198_/B _14176_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14177_/X
+ sky130_fd_sc_hd__o211a_1
X_11389_ hold5457/X _12338_/B _11388_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _11389_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13121_/X _13127_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17534_/D sky130_fd_sc_hd__o21a_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17936_ _17960_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13058_/X _16900_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
Xhold1009 hold1108/X vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__clkbuf_16
X_17867_ _17867_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16818_ _18019_/CLK _16818_/D vssd1 vssd1 vccd1 vccd1 _16818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17798_ _17869_/CLK _17798_/D vssd1 vssd1 vccd1 vccd1 _17798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16749_ _18014_/CLK _16749_/D vssd1 vssd1 vccd1 vccd1 _16749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ hold2186/X _09216_/B _09220_/X _12912_/A vssd1 vssd1 vccd1 vccd1 _09221_/X
+ sky130_fd_sc_hd__o211a_1
X_18419_ _18421_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _15535_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08103_ hold202/X hold238/X vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__nand2b_1
X_09083_ hold1123/X _09119_/A2 _09082_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08034_ hold2355/X _08033_/B _08033_/Y _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08034_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput70 input70/A vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 hold832/A vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 hold843/A vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 hold854/A vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/A vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/A vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold887 hold887/A vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold898 hold898/A vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _13070_/A _10025_/B _09984_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _16485_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2200 _08239_/X vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 _08091_/X vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08936_ _15374_/A hold640/X vssd1 vssd1 vccd1 vccd1 _16085_/D sky130_fd_sc_hd__and2_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2222 _09149_/X vssd1 vssd1 vccd1 vccd1 _16187_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2233 _17764_/Q vssd1 vssd1 vccd1 vccd1 hold2233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 _18063_/Q vssd1 vssd1 vccd1 vccd1 hold2244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 _14677_/X vssd1 vssd1 vccd1 vccd1 _18129_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2255 _09167_/X vssd1 vssd1 vccd1 vccd1 _16196_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1521 _16197_/Q vssd1 vssd1 vccd1 vccd1 hold1521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2266 _14269_/X vssd1 vssd1 vccd1 vccd1 _17933_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ _13037_/A hold444/X vssd1 vssd1 vccd1 vccd1 _16052_/D sky130_fd_sc_hd__and2_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1532 _18067_/Q vssd1 vssd1 vccd1 vccd1 hold1532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 _14049_/X vssd1 vssd1 vccd1 vccd1 _17828_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2288 _15873_/Q vssd1 vssd1 vccd1 vccd1 hold2288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 _08006_/X vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2299 _17991_/Q vssd1 vssd1 vccd1 vccd1 hold2299/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1554 _13922_/X vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1565 _18387_/Q vssd1 vssd1 vccd1 vccd1 hold1565/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1576 _08479_/X vssd1 vssd1 vccd1 vccd1 _15868_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ hold752/A hold764/A hold732/A hold689/A vssd1 vssd1 vccd1 vccd1 _14735_/A
+ sky130_fd_sc_hd__or4bb_4
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _12444_/A hold564/X vssd1 vssd1 vccd1 vccd1 _16018_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1587 _16200_/Q vssd1 vssd1 vccd1 vccd1 hold1587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1598 _08477_/X vssd1 vssd1 vccd1 vccd1 _15867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18438_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ hold1845/X hold5503/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_274_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18112_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09419_ _07804_/A hold5915/X _15304_/A _09418_/X vssd1 vssd1 vccd1 vccd1 _09419_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_203_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18350_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ hold2317/X hold4660/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10692_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _17308_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12361_ _13873_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _17277_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _15553_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14100_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11312_ hold1291/X hold3685/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__mux2_1
X_15080_ hold5981/X _15111_/B _15079_/X _15064_/A vssd1 vssd1 vccd1 vccd1 hold766/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12292_ hold5332/X _13798_/A2 _12291_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ hold2821/X _14040_/B _14030_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14031_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11243_ _18429_/Q hold3579/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ _16882_/Q _11177_/B _11204_/C vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__and3_1
XTAP_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4180 _11443_/X vssd1 vssd1 vccd1 vccd1 _16971_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10125_ _10533_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__or2_1
Xhold4191 _17203_/Q vssd1 vssd1 vccd1 vccd1 hold4191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _17293_/CLK _15982_/D vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
XTAP_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3490 _17714_/Q vssd1 vssd1 vccd1 vccd1 hold3490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17721_ _17721_/CLK _17721_/D vssd1 vssd1 vccd1 vccd1 _17721_/Q sky130_fd_sc_hd__dfxtp_1
X_10056_ _13262_/A _09960_/A _10055_/X vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__a21oi_1
X_14933_ hold3168/X _14952_/B _14932_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14933_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_21_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_21_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _17748_/CLK _17652_/D vssd1 vssd1 vccd1 vccd1 _17652_/Q sky130_fd_sc_hd__dfxtp_1
X_14864_ _14988_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _18223_/CLK _16603_/D vssd1 vssd1 vccd1 vccd1 _16603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ _17565_/Q _13800_/A _13814_/X vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__a21oi_1
X_14795_ hold1935/X _14826_/B _14794_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14795_/X
+ sky130_fd_sc_hd__o211a_1
X_17583_ _17711_/CLK _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16534_ _18186_/CLK _16534_/D vssd1 vssd1 vccd1 vccd1 _16534_/Q sky130_fd_sc_hd__dfxtp_1
X_13746_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__or2_1
X_10958_ hold2066/X hold3806/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _18376_/CLK _16465_/D vssd1 vssd1 vccd1 vccd1 _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _13746_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__or2_1
X_10889_ hold2413/X hold5042/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _18224_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _17317_/Q _09357_/A _09392_/A hold740/X vssd1 vssd1 vccd1 vccd1 _15416_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12628_ hold1100/X hold3340/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12628_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16396_ _18309_/CLK _16396_/D vssd1 vssd1 vccd1 vccd1 _16396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15347_ hold232/X _09357_/A _09386_/D hold258/X _15346_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/B sky130_fd_sc_hd__a221o_2
X_18135_ _18216_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ hold3100/X hold3599/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5809 hold5943/X vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__buf_1
XFILLER_0_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ hold539/X _15484_/A2 _09392_/D hold129/X vssd1 vssd1 vccd1 vccd1 _15278_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18066_ _18068_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
Xhold117 input10/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 input25/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14229_ hold1769/X _14216_/Y _14228_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _14229_/X
+ sky130_fd_sc_hd__o211a_1
X_17017_ _17767_/CLK _17017_/D vssd1 vssd1 vccd1 vccd1 _17017_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_78_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17499_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_60_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_60_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout608 _09361_/Y vssd1 vssd1 vccd1 vccd1 _15485_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_226_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout619 _09351_/Y vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09770_ hold2746/X _16414_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_225_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08721_ hold140/X hold193/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__mux2_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _18060_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08652_ _12404_/A hold835/X vssd1 vssd1 vccd1 vccd1 _15948_/D sky130_fd_sc_hd__and2_1
XFILLER_0_240_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08583_ _15264_/A hold231/X vssd1 vssd1 vccd1 vccd1 _15915_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09204_ _15533_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ hold2090/X _09177_/A2 _09134_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09066_ _15182_/A hold533/A vssd1 vssd1 vccd1 vccd1 _09066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08017_ _15531_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold640 hold640/A vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 hold651/A vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold673 hold673/A vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 hold684/A vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold695 hold695/A vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ hold1493/X _16480_/Q _10580_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__mux2_1
Xhold2030 _08459_/X vssd1 vssd1 vccd1 vccd1 _15858_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2041 _15544_/X vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08919_ _12416_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _16077_/D sky130_fd_sc_hd__and2_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2052 _08210_/X vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2063 _16206_/Q vssd1 vssd1 vccd1 vccd1 hold2063/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09899_ _18368_/Q hold3349/X _10019_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__mux2_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 _15723_/Q vssd1 vssd1 vccd1 vccd1 hold2074/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_232_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2085 _15795_/Q vssd1 vssd1 vccd1 vccd1 hold2085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1340 _15776_/Q vssd1 vssd1 vccd1 vccd1 hold1340/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1351 _07846_/X vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ hold2357/X hold5391/X _13862_/C vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__mux2_1
Xhold2096 _16182_/Q vssd1 vssd1 vccd1 vccd1 hold2096/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1362 _14051_/X vssd1 vssd1 vccd1 vccd1 _17829_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_455_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17721_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1373 _15589_/Q vssd1 vssd1 vccd1 vccd1 hold1373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _09415_/X vssd1 vssd1 vccd1 vccd1 _16293_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1395 _15797_/Q vssd1 vssd1 vccd1 vccd1 hold1395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ hold2864/X hold3724/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13600_ hold3519/X _13886_/B _13599_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13600_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10812_ _11115_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14580_ _15189_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11792_ _17088_/Q _11801_/B _11792_/C vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__and3_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13531_ hold5685/X _13829_/B _13530_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10743_ _11124_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _17413_/CLK _16250_/D vssd1 vssd1 vccd1 vccd1 _16250_/Q sky130_fd_sc_hd__dfxtp_1
X_13462_ hold4323/X _12374_/B _13461_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _13462_/X
+ sky130_fd_sc_hd__o211a_1
X_10674_ _11136_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15201_ _15201_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__or2_1
X_12413_ hold256/X hold780/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16181_ _17485_/CLK _16181_/D vssd1 vssd1 vccd1 vccd1 _16181_/Q sky130_fd_sc_hd__dfxtp_1
X_13393_ hold4449/X _13777_/A2 _13392_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15132_ hold1076/X _15167_/B _15131_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15132_/X
+ sky130_fd_sc_hd__o211a_1
X_12344_ _12344_/A _12344_/B _12344_/C vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15063_ _15225_/A hold1178/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15064_/B sky130_fd_sc_hd__mux2_1
X_12275_ hold2363/X hold4451/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14014_ _15521_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14014_/X sky130_fd_sc_hd__or2_1
X_11226_ hold4992/X _11670_/A _11225_/X vssd1 vssd1 vccd1 vccd1 _11226_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11157_ hold4911/X _11136_/A _11156_/X vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ hold5064/X _10625_/B _10107_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _17284_/CLK _15965_/D vssd1 vssd1 vccd1 vccd1 hold649/A sky130_fd_sc_hd__dfxtp_1
X_11088_ _11094_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__or2_1
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17704_ _17738_/CLK _17704_/D vssd1 vssd1 vccd1 vccd1 _17704_/Q sky130_fd_sc_hd__dfxtp_1
X_10039_ _10603_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _16503_/D sky130_fd_sc_hd__nor2_1
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14916_ _15185_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14916_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_196_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18356_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15896_ _17343_/CLK _15896_/D vssd1 vssd1 vccd1 vccd1 _15896_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17635_ _17667_/CLK _17635_/D vssd1 vssd1 vccd1 vccd1 _17635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_125_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14847_ hold1801/X _14880_/B _14846_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17566_ _17686_/CLK _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14778_ _15225_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16517_ _16517_/CLK _16517_/D vssd1 vssd1 vccd1 vccd1 _16517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13729_ hold5751/X _13832_/B _13728_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17497_ _17499_/CLK _17497_/D vssd1 vssd1 vccd1 vccd1 _17497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16448_ _18391_/CLK _16448_/D vssd1 vssd1 vccd1 vccd1 _16448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16379_ _18322_/CLK _16379_/D vssd1 vssd1 vccd1 vccd1 _16379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18118_ _18170_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5606 _11656_/X vssd1 vssd1 vccd1 vccd1 _17042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5617 _17238_/Q vssd1 vssd1 vccd1 vccd1 hold5617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5628 _11560_/X vssd1 vssd1 vccd1 vccd1 _17010_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5639 _17142_/Q vssd1 vssd1 vccd1 vccd1 hold5639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4905 _16921_/Q vssd1 vssd1 vccd1 vccd1 hold4905/X sky130_fd_sc_hd__dlygate4sd3_1
X_18049_ _18049_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4916 _12010_/X vssd1 vssd1 vccd1 vccd1 _17160_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4927 _17224_/Q vssd1 vssd1 vccd1 vccd1 hold4927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4938 _16625_/Q vssd1 vssd1 vccd1 vccd1 hold4938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4949 _10023_/Y vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 hold755/X vssd1 vssd1 vccd1 vccd1 _14326_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_240_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout416 _14107_/A2 vssd1 vssd1 vccd1 vccd1 _14094_/B sky130_fd_sc_hd__clkbuf_8
X_09822_ _09933_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__or2_1
Xfanout427 _13267_/S vssd1 vssd1 vccd1 vccd1 _13307_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout438 _13817_/C vssd1 vssd1 vccd1 vccd1 _13826_/C sky130_fd_sc_hd__buf_6
Xfanout449 _11150_/C vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__buf_6
XFILLER_0_226_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09753_ _11082_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09753_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08704_ _12438_/A hold403/X vssd1 vssd1 vccd1 vccd1 _15973_/D sky130_fd_sc_hd__and2_1
XFILLER_0_240_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09684_ _10470_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08635_ hold568/X hold617/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08636_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08566_ hold379/X hold694/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08497_ hold2439/X _08486_/B _08496_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08497_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09118_ _15559_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ hold3343/X _10598_/B _10389_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10390_/X
+ sky130_fd_sc_hd__o211a_1
X_09049_ _12430_/A hold579/X vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__and2_1
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12060_ _12231_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold470 hold470/A vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 hold492/A vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ hold5635/X _11201_/B _11010_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ hold3598/X _12961_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__mux2_1
X_15750_ _17701_/CLK _15750_/D vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _18203_/Q vssd1 vssd1 vccd1 vccd1 hold1170/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ hold3067/X _14720_/B _14700_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _14701_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 _16202_/Q vssd1 vssd1 vccd1 vccd1 hold1181/X sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _13716_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__or2_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 _15781_/Q vssd1 vssd1 vccd1 vccd1 hold1192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15681_ _17153_/CLK _15681_/D vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ hold3225/X _12892_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__mux2_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17420_/CLK _17420_/D vssd1 vssd1 vccd1 vccd1 _17420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14794_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__or2_1
X_11844_ _12219_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__or2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14563_ _14794_/A _14557_/Y hold1184/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14563_/X
+ sky130_fd_sc_hd__o211a_1
X_17351_ _17515_/CLK _17351_/D vssd1 vssd1 vccd1 vccd1 _17351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ hold3722/X _12057_/A _11774_/X vssd1 vssd1 vccd1 vccd1 _11775_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ _16320_/CLK hold826/X vssd1 vssd1 vccd1 vccd1 _16302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13514_ hold2999/X hold4171/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ hold4453/X _11753_/B _10725_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _10726_/X
+ sky130_fd_sc_hd__o211a_1
X_14494_ hold1640/X _14487_/B _14493_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _14494_/X
+ sky130_fd_sc_hd__o211a_1
X_17282_ _17607_/CLK _17282_/D vssd1 vssd1 vccd1 vccd1 _17282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ hold2158/X hold5695/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__mux2_1
X_16233_ _17413_/CLK _16233_/D vssd1 vssd1 vccd1 vccd1 _16233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ hold5483/X _11156_/B _10656_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ hold1575/X _17579_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__mux2_1
X_16164_ _18043_/CLK _16164_/D vssd1 vssd1 vccd1 vccd1 _16164_/Q sky130_fd_sc_hd__dfxtp_1
X_10588_ _18461_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _16686_/D sky130_fd_sc_hd__nor2_1
X_15115_ _15169_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15115_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12327_ hold3645/X _12231_/A _12326_/X vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__a21oi_1
X_16095_ _16095_/CLK _16095_/D vssd1 vssd1 vccd1 vccd1 hold660/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15046_ _15050_/A _15046_/B vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12258_ _13794_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11209_ _12340_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _16893_/D sky130_fd_sc_hd__nor2_1
X_12189_ _12285_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_377_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17728_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16997_ _17875_/CLK _16997_/D vssd1 vssd1 vccd1 vccd1 _16997_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_306_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17869_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _17298_/CLK _15948_/D vssd1 vssd1 vccd1 vccd1 hold834/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15879_ _17741_/CLK _15879_/D vssd1 vssd1 vccd1 vccd1 _15879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ hold2869/X _08440_/A2 _08419_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08420_/X
+ sky130_fd_sc_hd__o211a_1
X_17618_ _17650_/CLK _17618_/D vssd1 vssd1 vccd1 vccd1 _17618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__and2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17549_ _18215_/CLK _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08282_ hold752/A hold764/A hold732/X hold689/X vssd1 vssd1 vccd1 vccd1 hold733/A
+ sky130_fd_sc_hd__or4b_2
Xclkbuf_leaf_93_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18415_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17483_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5403 _16880_/Q vssd1 vssd1 vccd1 vccd1 hold5403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5414 _12094_/X vssd1 vssd1 vccd1 vccd1 _17188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5425 _16689_/Q vssd1 vssd1 vccd1 vccd1 hold5425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5436 _12067_/X vssd1 vssd1 vccd1 vccd1 _17179_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4702 _10620_/Y vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5447 _16831_/Q vssd1 vssd1 vccd1 vccd1 hold5447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4713 _16383_/Q vssd1 vssd1 vccd1 vccd1 hold4713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5458 _11389_/X vssd1 vssd1 vccd1 vccd1 _16953_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4724 _09691_/X vssd1 vssd1 vccd1 vccd1 _16387_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5469 _17085_/Q vssd1 vssd1 vccd1 vccd1 hold5469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4735 _16378_/Q vssd1 vssd1 vccd1 vccd1 hold4735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4746 _10480_/X vssd1 vssd1 vccd1 vccd1 _16650_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4757 _16616_/Q vssd1 vssd1 vccd1 vccd1 hold4757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4768 _09673_/X vssd1 vssd1 vccd1 vccd1 _16381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4779 _17116_/Q vssd1 vssd1 vccd1 vccd1 hold4779/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout202 _11584_/A2 vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__clkbuf_8
Xfanout213 _10004_/B vssd1 vssd1 vccd1 vccd1 _10034_/B sky130_fd_sc_hd__buf_4
Xfanout224 _10468_/A2 vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout235 _10037_/B vssd1 vssd1 vccd1 vccd1 _10565_/B sky130_fd_sc_hd__buf_4
Xfanout246 _09494_/X vssd1 vssd1 vccd1 vccd1 fanout246/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09805_ hold3349/X _10013_/B _09804_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09805_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout257 _13623_/A vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__buf_2
Xfanout268 _11070_/A vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__buf_4
Xfanout279 fanout334/X vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__buf_4
X_07997_ hold915/X _08045_/B vssd1 vssd1 vccd1 vccd1 _07997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09736_ hold4535/X _09832_/A2 _09735_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09736_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ hold3635/X _10049_/B _09666_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09667_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08618_ _09015_/A hold185/X vssd1 vssd1 vccd1 vccd1 _15931_/D sky130_fd_sc_hd__and2_1
XFILLER_0_194_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ hold4123/X _10004_/B _09597_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09598_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08549_ _12436_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _15898_/D sky130_fd_sc_hd__and2_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ hold5627/X _11753_/B _11559_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11560_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ hold1977/X _16661_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ hold5266/X _12317_/B _11490_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11491_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ _13230_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__or2_1
X_10442_ hold1094/X _16638_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ _13161_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__and2_1
XFILLER_0_165_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ hold3114/X _16615_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ hold4940/X _13811_/B _12111_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _12112_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5970 _13040_/X vssd1 vssd1 vccd1 vccd1 hold931/A sky130_fd_sc_hd__dlygate4sd3_1
X_13092_ hold3679/X _13091_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_2
Xhold5981 _18322_/Q vssd1 vssd1 vccd1 vccd1 hold5981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5992 _17941_/Q vssd1 vssd1 vccd1 vccd1 hold5992/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12043_ hold4191/X _13871_/B _12042_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12043_/X
+ sky130_fd_sc_hd__o211a_1
X_16920_ _17869_/CLK _16920_/D vssd1 vssd1 vccd1 vccd1 _16920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ _18052_/CLK _16851_/D vssd1 vssd1 vccd1 vccd1 _16851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 _08147_/A vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15802_ _17745_/CLK _15802_/D vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout791 _13935_/A vssd1 vssd1 vccd1 vccd1 _14203_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16782_ _18060_/CLK _16782_/D vssd1 vssd1 vccd1 vccd1 _16782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13994_ _14782_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15733_ _17736_/CLK _15733_/D vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12999_/A _12945_/B vssd1 vssd1 vccd1 vccd1 _17491_/D sky130_fd_sc_hd__and2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18452_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _17872_/CLK _15664_/D vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12990_/A _12876_/B vssd1 vssd1 vccd1 vccd1 _17468_/D sky130_fd_sc_hd__and2_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17403_ _18453_/CLK _17403_/D vssd1 vssd1 vccd1 vccd1 _17403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14615_ hold2246/X _14610_/B _14614_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14615_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18383_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
X_11827_ hold5072/X _12308_/B _11826_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11827_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _17718_/CLK _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ _17334_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 _17334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14546_ hold1532/X _14541_/B _14545_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14546_/X
+ sky130_fd_sc_hd__o211a_1
X_11758_ _12340_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _17076_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_126_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ hold2974/X hold4670/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__mux2_1
X_17265_ _17265_/CLK _17265_/D vssd1 vssd1 vccd1 vccd1 _17265_/Q sky130_fd_sc_hd__dfxtp_1
X_11689_ hold5469/X _12329_/B _11688_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11689_/X
+ sky130_fd_sc_hd__o211a_1
X_14477_ _15103_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14477_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ _17878_/CLK _16216_/D vssd1 vssd1 vccd1 vccd1 _16216_/Q sky130_fd_sc_hd__dfxtp_1
X_13428_ _13713_/A _13428_/B vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or2_1
X_17196_ _17253_/CLK _17196_/D vssd1 vssd1 vccd1 vccd1 _17196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16147_ _17343_/CLK _16147_/D vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13359_ _13761_/A _13359_/B vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4009 _10546_/X vssd1 vssd1 vccd1 vccd1 _16672_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16078_ _18415_/CLK _16078_/D vssd1 vssd1 vccd1 vccd1 _16078_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3308 _17438_/Q vssd1 vssd1 vccd1 vccd1 hold3308/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3319 _17462_/Q vssd1 vssd1 vccd1 vccd1 hold3319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07920_ _15543_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07920_/Y sky130_fd_sc_hd__nand2_1
X_15029_ _15191_/A hold2146/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15030_/B sky130_fd_sc_hd__mux2_1
Xhold2607 _15580_/Q vssd1 vssd1 vccd1 vccd1 hold2607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 _17905_/Q vssd1 vssd1 vccd1 vccd1 hold2618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _15120_/X vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1906 _18242_/Q vssd1 vssd1 vccd1 vccd1 hold1906/X sky130_fd_sc_hd__dlygate4sd3_1
X_07851_ _15529_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07851_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_140_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18364_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1917 _15683_/Q vssd1 vssd1 vccd1 vccd1 hold1917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 _14655_/X vssd1 vssd1 vccd1 vccd1 _18118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _17909_/Q vssd1 vssd1 vccd1 vccd1 hold1939/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput2 input2/A vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07782_ hold246/X vssd1 vssd1 vccd1 vccd1 _07782_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ hold1906/X _13118_/A _10001_/C vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09452_ _09456_/C _09456_/D _09456_/B vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_189_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _15517_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09383_ _15480_/A _09383_/B _09383_/C _09383_/D vssd1 vssd1 vccd1 vccd1 _09383_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_231_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ hold1559/X _08323_/B _08333_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08265_ hold2000/X _08268_/B _08264_/Y _08351_/A vssd1 vssd1 vccd1 vccd1 _08265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ hold2945/X _08213_/B _08195_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5200 _16942_/Q vssd1 vssd1 vccd1 vccd1 hold5200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5211 _10273_/X vssd1 vssd1 vccd1 vccd1 _16581_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5222 _17006_/Q vssd1 vssd1 vccd1 vccd1 hold5222/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5233 _11812_/X vssd1 vssd1 vccd1 vccd1 _17094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_299_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5244 _16646_/Q vssd1 vssd1 vccd1 vccd1 hold5244/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5255 _11935_/X vssd1 vssd1 vccd1 vccd1 _17135_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4510 _10729_/X vssd1 vssd1 vccd1 vccd1 _16733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4521 _17640_/Q vssd1 vssd1 vccd1 vccd1 hold4521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5266 _17019_/Q vssd1 vssd1 vccd1 vccd1 hold5266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5277 _10900_/X vssd1 vssd1 vccd1 vccd1 _16790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4532 _11029_/X vssd1 vssd1 vccd1 vccd1 _16833_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_228_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18131_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_219_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5288 _16324_/Q vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4543 _17144_/Q vssd1 vssd1 vccd1 vccd1 hold4543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4554 _10936_/X vssd1 vssd1 vccd1 vccd1 _16802_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3820 _09862_/X vssd1 vssd1 vccd1 vccd1 _16444_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5299 _13318_/X vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4565 _17742_/Q vssd1 vssd1 vccd1 vccd1 hold4565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4576 _13573_/X vssd1 vssd1 vccd1 vccd1 _17644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3831 _16933_/Q vssd1 vssd1 vccd1 vccd1 hold3831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4587 hold5871/X vssd1 vssd1 vccd1 vccd1 hold5872/A sky130_fd_sc_hd__buf_4
Xhold3842 _10897_/X vssd1 vssd1 vccd1 vccd1 _16789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4598 _10032_/Y vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3853 _11799_/Y vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3864 _16501_/Q vssd1 vssd1 vccd1 vccd1 _10031_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3875 _10261_/X vssd1 vssd1 vccd1 vccd1 _16577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3886 _16494_/Q vssd1 vssd1 vccd1 vccd1 hold3886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3897 _15333_/X vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ hold3038/X hold3405/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__mux2_1
X_10991_ hold1901/X hold3841/X _11093_/S vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ hold1196/X _17421_/Q _12748_/S vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__mux2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ hold2188/X _17398_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ hold1998/X _14446_/A2 _14399_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14400_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ hold2023/X _17028_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ hold893/X _09367_/A _09392_/A hold804/X vssd1 vssd1 vccd1 vccd1 _15380_/X
+ sky130_fd_sc_hd__a22o_1
X_12592_ hold2457/X _17375_/Q _12967_/S vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14331_ hold1458/X _14326_/B _14330_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14331_/X
+ sky130_fd_sc_hd__o211a_1
X_11543_ hold2271/X hold5292/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14262_ _15103_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or2_1
X_17050_ _17896_/CLK _17050_/D vssd1 vssd1 vccd1 vccd1 _17050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11474_ hold2276/X _16982_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13213_ _13212_/X hold3549/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__mux2_2
X_16001_ _18406_/CLK _16001_/D vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__dfxtp_1
X_10425_ _10830_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ hold2735/X _14198_/B _14192_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13144_ _13137_/X _13143_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17536_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _10998_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13074_/X _16902_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__mux2_1
X_17952_ _17952_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
X_10287_ _11097_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12026_ hold2648/X _17166_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__mux2_1
X_16903_ _17814_/CLK _16903_/D vssd1 vssd1 vccd1 vccd1 _16903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17883_ _17883_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16834_ _18035_/CLK _16834_/D vssd1 vssd1 vccd1 vccd1 _16834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16765_ _17966_/CLK _16765_/D vssd1 vssd1 vccd1 vccd1 _16765_/Q sky130_fd_sc_hd__dfxtp_1
X_13977_ hold1873/X _13986_/B _13976_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _13977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ _17188_/CLK _15716_/D vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12928_ hold1026/X hold3251/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_220_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16696_ _17968_/CLK _16696_/D vssd1 vssd1 vccd1 vccd1 _16696_/Q sky130_fd_sc_hd__dfxtp_1
X_18435_ _18435_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
X_15647_ _17194_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ hold2090/X hold3297/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ _18366_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15578_ _17742_/CLK _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _17320_/CLK hold102/X vssd1 vssd1 vccd1 vccd1 _17317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14529_ _14529_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14529_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18297_ _18391_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _15509_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__or2_1
X_17248_ _17280_/CLK _17248_/D vssd1 vssd1 vccd1 vccd1 _17248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17179_ _17179_/CLK _17179_/D vssd1 vssd1 vccd1 vccd1 _17179_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_392_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17895_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_321_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17870_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3105 _14532_/X vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3116 _18141_/Q vssd1 vssd1 vccd1 vccd1 hold3116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3127 _10026_/Y vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ _15414_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _16093_/D sky130_fd_sc_hd__and2_1
Xhold3138 _17504_/Q vssd1 vssd1 vccd1 vccd1 hold3138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2404 _07973_/X vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 _17468_/Q vssd1 vssd1 vccd1 vccd1 hold3149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _14025_/X vssd1 vssd1 vccd1 vccd1 _17816_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07903_ hold2793/X _07924_/B _07902_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07903_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2426 _17821_/Q vssd1 vssd1 vccd1 vccd1 hold2426/X sky130_fd_sc_hd__dlygate4sd3_1
X_08883_ _15264_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _16059_/D sky130_fd_sc_hd__and2_1
Xhold2437 _08198_/X vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 _14963_/X vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _14613_/X vssd1 vssd1 vccd1 vccd1 _18098_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2459 _15642_/Q vssd1 vssd1 vccd1 vccd1 hold2459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _16201_/Q vssd1 vssd1 vccd1 vccd1 hold1714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 hold1725/A vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__buf_12
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07834_ hold1444/X _07865_/B _07833_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _07834_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1736 _08487_/X vssd1 vssd1 vccd1 vccd1 _15872_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 _07937_/X vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1758 _14623_/X vssd1 vssd1 vccd1 vccd1 _18103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _17914_/Q vssd1 vssd1 vccd1 vccd1 hold1769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_154_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09504_ _09984_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _07785_/Y hold850/X _15344_/A _09434_/X vssd1 vssd1 vccd1 vccd1 hold851/A
+ sky130_fd_sc_hd__o211a_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_164_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _15541_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _15519_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__or2_1
XANTENNA_40 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _14862_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__or2_1
XANTENNA_73 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 hold181/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_409_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17821_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_95 hold1152/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08179_ _15513_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5030 _17724_/Q vssd1 vssd1 vccd1 vccd1 hold5030/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5041 _09796_/X vssd1 vssd1 vccd1 vccd1 _16422_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10210_ hold3742/X _10628_/B _10209_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5052 _16368_/Q vssd1 vssd1 vccd1 vccd1 hold5052/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ hold4670/X _11121_/A _11189_/X vssd1 vssd1 vccd1 vccd1 _11190_/Y sky130_fd_sc_hd__a21oi_1
Xhold5063 _11434_/X vssd1 vssd1 vccd1 vccd1 _16968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5074 _17084_/Q vssd1 vssd1 vccd1 vccd1 hold5074/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5085 _11077_/X vssd1 vssd1 vccd1 vccd1 _16849_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4340 _17152_/Q vssd1 vssd1 vccd1 vccd1 hold4340/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10141_ hold5433/X _10619_/B _10140_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5096 _17227_/Q vssd1 vssd1 vccd1 vccd1 hold5096/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4351 _11581_/X vssd1 vssd1 vccd1 vccd1 _17017_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4362 _16871_/Q vssd1 vssd1 vccd1 vccd1 hold4362/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4373 _13594_/X vssd1 vssd1 vccd1 vccd1 _17651_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4384 _17733_/Q vssd1 vssd1 vccd1 vccd1 hold4384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3650 _13860_/Y vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4395 _17670_/Q vssd1 vssd1 vccd1 vccd1 hold4395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10072_ _11194_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _16514_/D sky130_fd_sc_hd__nor2_1
Xhold3661 _17395_/Q vssd1 vssd1 vccd1 vccd1 hold3661/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3672 _16439_/Q vssd1 vssd1 vccd1 vccd1 hold3672/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3683 _17123_/Q vssd1 vssd1 vccd1 vccd1 hold3683/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3694 _12719_/X vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_11_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_11_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_13900_ _15189_/A hold3014/X hold124/X vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__mux2_1
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2960 _15530_/X vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14880_ _15004_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__nand2_1
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2971 _18095_/Q vssd1 vssd1 vccd1 vccd1 hold2971/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2982 _14965_/X vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2993 _16266_/Q vssd1 vssd1 vccd1 vccd1 hold2993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13831_ _13864_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _17730_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_216_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16550_ _18170_/CLK _16550_/D vssd1 vssd1 vccd1 vccd1 _16550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _11070_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__or2_1
X_13762_ hold4479/X _13856_/B _13761_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15517_/A hold1949/X hold691/X vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ hold3696/X _12712_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__mux2_1
X_16481_ _16517_/CLK _16481_/D vssd1 vssd1 vccd1 vccd1 _16481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ hold4197/X _13883_/B _13692_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _18220_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15432_ _15480_/A _15432_/B _15432_/C _15432_/D vssd1 vssd1 vccd1 vccd1 _15432_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ hold3527/X _12643_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18151_ _18175_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_15363_ _15490_/A1 _15355_/X _15362_/X _15490_/B1 hold5870/A vssd1 vssd1 vccd1 vccd1
+ _15363_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12575_ hold3585/X _12574_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17102_ _17166_/CLK _17102_/D vssd1 vssd1 vccd1 vccd1 _17102_/Q sky130_fd_sc_hd__dfxtp_1
X_14314_ _14529_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14314_/X sky130_fd_sc_hd__or2_1
X_18082_ _18224_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _12204_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__or2_1
X_15294_ _15374_/A _15294_/B vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__and2_1
XFILLER_0_123_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _17815_/CLK _17033_/D vssd1 vssd1 vccd1 vccd1 _17033_/Q sky130_fd_sc_hd__dfxtp_1
X_14245_ hold2636/X _14266_/B _14244_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14245_/X
+ sky130_fd_sc_hd__o211a_1
X_11457_ _11553_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ hold4849/X _11192_/B _10407_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10408_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_50_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_50_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14176_ _14246_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14176_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ _12243_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ hold4829/X _10477_/A2 _10338_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10339_/X
+ sky130_fd_sc_hd__o211a_1
X_13127_ _13199_/A1 _13125_/X _13126_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _17558_/Q _17092_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__mux2_1
X_17935_ _17935_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12009_ _13716_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__or2_1
X_17866_ _17898_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ _18050_/CLK _16817_/D vssd1 vssd1 vccd1 vccd1 _16817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17797_ _17891_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16748_ _18305_/CLK _16748_/D vssd1 vssd1 vccd1 vccd1 _16748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16679_ _18296_/CLK _16679_/D vssd1 vssd1 vccd1 vccd1 _16679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _15549_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__or2_1
X_18418_ _18418_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09151_ hold2806/X _09164_/B _09150_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _09151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18349_ _18349_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08102_ hold689/A hold764/A hold732/A hold752/A vssd1 vssd1 vccd1 vccd1 hold238/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _15523_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08033_ _14774_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08033_/Y sky130_fd_sc_hd__nand2_1
Xhold800 hold800/A vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_6
Xhold811 hold811/A vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput71 wb_rst_i vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold822 slv_done vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 hold844/A vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/A vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 hold866/A vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold877 hold877/A vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 hold888/A vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__or2_1
Xhold899 hold899/A vssd1 vssd1 vccd1 vccd1 hold899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2201 _15593_/Q vssd1 vssd1 vccd1 vccd1 hold2201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2212 _15577_/Q vssd1 vssd1 vccd1 vccd1 hold2212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ hold554/X hold639/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold640/A sky130_fd_sc_hd__mux2_1
Xhold2223 _15733_/Q vssd1 vssd1 vccd1 vccd1 hold2223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2234 _18336_/Q vssd1 vssd1 vccd1 vccd1 hold2234/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1500 _15536_/X vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 _14538_/X vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2256 _15633_/Q vssd1 vssd1 vccd1 vccd1 hold2256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 _17955_/Q vssd1 vssd1 vccd1 vccd1 hold1511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2267 _15676_/Q vssd1 vssd1 vccd1 vccd1 hold2267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _09169_/X vssd1 vssd1 vccd1 vccd1 _16197_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ hold150/X hold443/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold444/A sky130_fd_sc_hd__mux2_1
Xhold1533 _14546_/X vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 _17876_/Q vssd1 vssd1 vccd1 vccd1 hold2278/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1544 _18426_/Q vssd1 vssd1 vccd1 vccd1 hold1544/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2289 _08489_/X vssd1 vssd1 vccd1 vccd1 _15873_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 _18181_/Q vssd1 vssd1 vccd1 vccd1 hold1555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1566 _15214_/X vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07817_ _07817_/A _07817_/B _07817_/C _07817_/D vssd1 vssd1 vccd1 vccd1 _09366_/A
+ sky130_fd_sc_hd__or4_4
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08797_ hold554/X hold563/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold564/A sky130_fd_sc_hd__mux2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1577 _15783_/Q vssd1 vssd1 vccd1 vccd1 hold1577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1588 _09175_/X vssd1 vssd1 vccd1 vccd1 _16200_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 _18254_/Q vssd1 vssd1 vccd1 vccd1 hold1599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _09438_/B _09418_/B vssd1 vssd1 vccd1 vccd1 _09418_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10690_ hold5429/X _11168_/B _10689_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _10690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _09366_/A _09351_/B _09364_/B vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_30_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ hold3625/X _13773_/A _12359_/X vssd1 vssd1 vccd1 vccd1 _12360_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_243_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ hold4354/X _11584_/A2 _11310_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ _13797_/A _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__or2_1
X_14030_ _15537_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14030_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11242_ hold3928/X _11617_/A2 _11241_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11242_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11173_ _12310_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _16881_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_219_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4170 _10264_/X vssd1 vssd1 vccd1 vccd1 _16578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4181 _16427_/Q vssd1 vssd1 vccd1 vccd1 hold4181/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10124_ hold3189/X hold4630/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__mux2_1
XTAP_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4192 _12043_/X vssd1 vssd1 vccd1 vccd1 _17171_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15981_ _16128_/CLK _15981_/D vssd1 vssd1 vccd1 vccd1 hold714/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _17725_/CLK _17720_/D vssd1 vssd1 vccd1 vccd1 _17720_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3480 _17219_/Q vssd1 vssd1 vccd1 vccd1 hold3480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ _16509_/Q _10055_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__and3_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _15201_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__or2_1
Xhold3491 _13687_/X vssd1 vssd1 vccd1 vccd1 _17682_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _17683_/CLK _17651_/D vssd1 vssd1 vccd1 vccd1 _17651_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2790 _09227_/X vssd1 vssd1 vccd1 vccd1 _16225_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ hold2546/X _14882_/B _14862_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14863_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ _18216_/CLK _16602_/D vssd1 vssd1 vccd1 vccd1 _16602_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13814_ _13814_/A _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13814_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17582_ _17742_/CLK _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
X_14794_ _14794_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _18193_/CLK _16533_/D vssd1 vssd1 vccd1 vccd1 _16533_/Q sky130_fd_sc_hd__dfxtp_1
X_13745_ hold1130/X _17702_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__mux2_1
X_10957_ hold4299/X _11147_/B _10956_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ _18363_/CLK _16464_/D vssd1 vssd1 vccd1 vccd1 _16464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13676_ _15760_/Q _17679_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ hold5523/X _11210_/B _10887_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__o211a_1
X_18203_ _18205_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
X_15415_ hold385/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _12789_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _17385_/D sky130_fd_sc_hd__and2_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _18370_/CLK _16395_/D vssd1 vssd1 vccd1 vccd1 _16395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _18180_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
X_15346_ _17338_/Q _15448_/B1 _09362_/D _16115_/Q vssd1 vssd1 vccd1 vccd1 _15346_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12558_ _12960_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _17362_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18065_ _18065_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
X_11509_ hold4319/X _12365_/B _11508_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11509_/X
+ sky130_fd_sc_hd__o211a_1
X_15277_ hold475/X _15487_/A2 _15484_/B1 _17311_/Q _15276_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ hold50/X _12509_/A2 _12507_/A3 _12488_/X _09055_/A vssd1 vssd1 vccd1 vccd1
+ hold51/A sky130_fd_sc_hd__o311a_1
Xhold107 hold178/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 hold38/X vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__buf_4
XFILLER_0_145_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _17862_/CLK _17016_/D vssd1 vssd1 vccd1 vccd1 _17016_/Q sky130_fd_sc_hd__dfxtp_1
X_14228_ _15519_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ hold1861/X _14148_/B _14158_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14159_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout609 _09361_/Y vssd1 vssd1 vccd1 vccd1 _09362_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08720_ _12418_/A hold715/X vssd1 vssd1 vccd1 vccd1 _15981_/D sky130_fd_sc_hd__and2_1
X_17918_ _18337_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_241_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08651_ hold210/X hold834/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold835/A sky130_fd_sc_hd__mux2_1
X_17849_ _17975_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08582_ hold222/X hold230/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ hold2242/X _09218_/B _09202_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09203_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09134_ _15517_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _14555_/C hold532/X vssd1 vssd1 vccd1 vccd1 hold533/A sky130_fd_sc_hd__or2_4
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08016_ hold2785/X _08029_/B _08015_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _08016_/X
+ sky130_fd_sc_hd__o211a_1
Xhold630 hold630/A vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 hold652/A vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/A vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold685 hold685/A vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09967_ hold3621/X _10601_/B _09966_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09967_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2020 _15822_/Q vssd1 vssd1 vccd1 vccd1 hold2020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 _17822_/Q vssd1 vssd1 vccd1 vccd1 hold2031/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2042 _15617_/Q vssd1 vssd1 vccd1 vccd1 hold2042/X sky130_fd_sc_hd__dlygate4sd3_1
X_08918_ hold578/X hold627/X _08928_/S vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__mux2_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 _15806_/Q vssd1 vssd1 vccd1 vccd1 hold2053/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09898_ hold3363/X _10013_/B _09897_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _09898_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _09189_/X vssd1 vssd1 vccd1 vccd1 _16206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1330 _09405_/X vssd1 vssd1 vccd1 vccd1 _16288_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 _18037_/Q vssd1 vssd1 vccd1 vccd1 hold2075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2086 _08324_/X vssd1 vssd1 vccd1 vccd1 _15795_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _08286_/X vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 _15804_/Q vssd1 vssd1 vccd1 vccd1 hold1352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 _09139_/X vssd1 vssd1 vccd1 vccd1 _16182_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08849_ _12412_/A hold902/X vssd1 vssd1 vccd1 vccd1 _16043_/D sky130_fd_sc_hd__and2_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1363 _15678_/Q vssd1 vssd1 vccd1 vccd1 hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _07891_/X vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _16173_/Q vssd1 vssd1 vccd1 vccd1 hold1385/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1396 _08328_/X vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ hold5639/X _12052_/A2 _11859_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11860_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ hold2092/X hold4403/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__mux2_1
X_11791_ _12367_/A _11791_/B vssd1 vssd1 vccd1 vccd1 _17087_/D sky130_fd_sc_hd__nor2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _13734_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10742_ hold2387/X hold4919/X _11768_/C vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_424_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17188_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10673_ hold1593/X hold4903/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__mux2_1
X_13461_ _13461_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13461_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ hold1983/X _15219_/B _15199_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15200_/X
+ sky130_fd_sc_hd__o211a_1
X_12412_ _12412_/A hold796/X vssd1 vssd1 vccd1 vccd1 _17299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16180_ _17485_/CLK _16180_/D vssd1 vssd1 vccd1 vccd1 _16180_/Q sky130_fd_sc_hd__dfxtp_1
X_13392_ _13761_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15131_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15131_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12343_ _12367_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _17271_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15062_ _15062_/A _15062_/B vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ hold3496/X _12274_/A2 _12273_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12274_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11225_ _16899_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__and3_1
X_14013_ hold1210/X _14040_/B _14012_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _14013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11156_ _16876_/Q _11156_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__and3_1
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10107_ _10533_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15964_ _16131_/CLK _15964_/D vssd1 vssd1 vccd1 vccd1 hold781/A sky130_fd_sc_hd__dfxtp_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ hold3120/X _16853_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__mux2_1
XTAP_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17703_/CLK _17703_/D vssd1 vssd1 vccd1 vccd1 _17703_/Q sky130_fd_sc_hd__dfxtp_1
X_10038_ _13214_/A _09960_/A _10037_/X vssd1 vssd1 vccd1 vccd1 _10038_/Y sky130_fd_sc_hd__a21oi_1
X_14915_ hold1906/X _14946_/B _14914_/X _14915_/C1 vssd1 vssd1 vccd1 vccd1 _14915_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15895_ _17346_/CLK _15895_/D vssd1 vssd1 vccd1 vccd1 _15895_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _17666_/CLK _17634_/D vssd1 vssd1 vccd1 vccd1 _17634_/Q sky130_fd_sc_hd__dfxtp_1
X_14846_ _15131_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__or2_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17565_ _17725_/CLK _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
X_14777_ hold2516/X _14772_/B _14776_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14777_/X
+ sky130_fd_sc_hd__o211a_1
X_11989_ hold4401/X _13877_/B _11988_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _18234_/CLK _16516_/D vssd1 vssd1 vccd1 vccd1 _16516_/Q sky130_fd_sc_hd__dfxtp_1
X_13728_ _13767_/A _13728_/B vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__or2_1
X_17496_ _17496_/CLK _17496_/D vssd1 vssd1 vccd1 vccd1 _17496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_165_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18371_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16447_ _18294_/CLK _16447_/D vssd1 vssd1 vccd1 vccd1 _16447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13659_ _13791_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16378_ _18353_/CLK _16378_/D vssd1 vssd1 vccd1 vccd1 _16378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18117_ _18159_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15329_ hold418/X _15485_/A2 _15488_/A2 hold387/X _15328_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5607 _16803_/Q vssd1 vssd1 vccd1 vccd1 hold5607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5618 _12148_/X vssd1 vssd1 vccd1 vccd1 _17206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5629 _17080_/Q vssd1 vssd1 vccd1 vccd1 hold5629/X sky130_fd_sc_hd__dlygate4sd3_1
X_18048_ _18050_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4906 _11772_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4917 _17194_/Q vssd1 vssd1 vccd1 vccd1 hold4917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4928 _12106_/X vssd1 vssd1 vccd1 vccd1 _17192_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4939 _10309_/X vssd1 vssd1 vccd1 vccd1 _16593_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout406 _14280_/B vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__buf_6
XFILLER_0_201_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ hold2628/X _16431_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__mux2_1
Xfanout417 _14054_/Y vssd1 vssd1 vccd1 vccd1 _14107_/A2 sky130_fd_sc_hd__buf_6
Xfanout428 _13054_/X vssd1 vssd1 vccd1 vccd1 _13181_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout439 _13817_/C vssd1 vssd1 vccd1 vccd1 _13832_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09752_ hold2973/X hold4819/X _11177_/C vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08703_ hold402/X _15973_/Q _08721_/S vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09683_ _18296_/Q hold3708/X _10571_/C vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _12531_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _15939_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _15491_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _15906_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08496_ _14782_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09117_ hold1385/X _09119_/A2 _09116_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09048_ hold578/X _16141_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold471 hold471/A vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 hold482/A vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _11106_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout940 _15205_/A vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__buf_8
XFILLER_0_239_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12961_ hold2991/X hold3289/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__mux2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _07929_/X vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1171 _14831_/X vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ _15201_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14700_/X sky130_fd_sc_hd__or2_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 _09181_/X vssd1 vssd1 vccd1 vccd1 _16202_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ hold2601/X _17128_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__mux2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _17245_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _08296_/X vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ hold2739/X _17475_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14631_ hold1789/X _14666_/B _14630_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14631_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11843_ hold2118/X hold4871/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17350_ _18398_/CLK _17350_/D vssd1 vssd1 vccd1 vccd1 _17350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ hold690/X _14573_/B hold1183/X vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__a21o_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _17082_/Q _12344_/B _12344_/C vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16320_/CLK hold821/X vssd1 vssd1 vccd1 vccd1 _16301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ hold4083/X _13814_/B _13512_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _13513_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17281_ _17585_/CLK _17281_/D vssd1 vssd1 vccd1 vccd1 _17281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _11115_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__or2_1
X_14493_ _15173_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14493_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16232_ _17413_/CLK _16232_/D vssd1 vssd1 vccd1 vccd1 _16232_/Q sky130_fd_sc_hd__dfxtp_1
X_13444_ hold5745/X _13832_/B _13443_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10656_ _11136_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _17499_/CLK _16163_/D vssd1 vssd1 vccd1 vccd1 _16163_/Q sky130_fd_sc_hd__dfxtp_1
X_10587_ hold4687/X _10533_/A _10586_/X vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13375_ hold3504/X _13886_/B _13374_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15114_ hold1102/X _15113_/B _15113_/Y _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15114_/X
+ sky130_fd_sc_hd__o211a_1
X_12326_ _17266_/Q _12347_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__and3_1
X_16094_ _16127_/CLK _16094_/D vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15045_ _15099_/A hold2898/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15046_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_239_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ hold2872/X _17243_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ hold4962/X _11694_/A _11207_/X vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__a21oi_1
X_12188_ hold2021/X _17220_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11139_ _11139_/A _11139_/B vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__or2_1
X_16996_ _17842_/CLK _16996_/D vssd1 vssd1 vccd1 vccd1 _16996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ _18402_/CLK _15947_/D vssd1 vssd1 vccd1 vccd1 hold643/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _17650_/CLK _15878_/D vssd1 vssd1 vccd1 vccd1 _15878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_346_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_231_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14829_ hold1607/X _14828_/B _14828_/Y _14829_/C1 vssd1 vssd1 vccd1 vccd1 _14829_/X
+ sky130_fd_sc_hd__o211a_1
X_17617_ _17650_/CLK _17617_/D vssd1 vssd1 vccd1 vccd1 _17617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08350_ _14854_/A hold1059/X hold134/X vssd1 vssd1 vccd1 vccd1 _08350_/X sky130_fd_sc_hd__mux2_1
X_17548_ _18215_/CLK _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ hold1793/X _08268_/B _08280_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _08281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ _17479_/CLK _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5404 _11074_/X vssd1 vssd1 vccd1 vccd1 _16848_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5415 _16749_/Q vssd1 vssd1 vccd1 vccd1 hold5415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5426 _10501_/X vssd1 vssd1 vccd1 vccd1 _16657_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5437 _17014_/Q vssd1 vssd1 vccd1 vccd1 hold5437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4703 _16851_/Q vssd1 vssd1 vccd1 vccd1 hold4703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5448 _10927_/X vssd1 vssd1 vccd1 vccd1 _16799_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4714 _09583_/X vssd1 vssd1 vccd1 vccd1 _16351_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5459 _17622_/Q vssd1 vssd1 vccd1 vccd1 hold5459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4725 _16529_/Q vssd1 vssd1 vccd1 vccd1 hold4725/X sky130_fd_sc_hd__buf_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4736 _09568_/X vssd1 vssd1 vccd1 vccd1 _16346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_62_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18038_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4747 _17581_/Q vssd1 vssd1 vccd1 vccd1 hold4747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4758 _10282_/X vssd1 vssd1 vccd1 vccd1 _16584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4769 _16387_/Q vssd1 vssd1 vccd1 vccd1 hold4769/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout203 _11584_/A2 vssd1 vssd1 vccd1 vccd1 _11801_/B sky130_fd_sc_hd__buf_2
Xfanout214 _09832_/A2 vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout225 _10468_/A2 vssd1 vssd1 vccd1 vccd1 _10598_/B sky130_fd_sc_hd__buf_4
Xfanout236 _10037_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__buf_4
XFILLER_0_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09804_ _09918_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__or2_1
Xfanout247 _13800_/A vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout258 fanout334/X vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__buf_4
Xfanout269 _11139_/A vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07996_ hold1767/X _08029_/B _07995_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _07996_/X
+ sky130_fd_sc_hd__o211a_1
X_09735_ _09843_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__or2_1
XFILLER_0_236_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _09954_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08617_ hold163/X hold184/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09987_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08548_ hold174/X hold234/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08479_ hold1575/X _08488_/B _08478_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08479_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ hold4813/X _10649_/B _10509_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _12285_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ hold5098/X _10631_/B _10440_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _13153_/X _13159_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17538_/D sky130_fd_sc_hd__o21a_1
X_10372_ hold5244/X _10468_/A2 _10371_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _10372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ _13716_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__or2_1
Xhold5960 data_in[17] vssd1 vssd1 vccd1 vccd1 hold376/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13091_ _13090_/X _16904_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
Xhold5971 data_in[26] vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5982 _18292_/Q vssd1 vssd1 vccd1 vccd1 hold5982/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5993 _18341_/Q vssd1 vssd1 vccd1 vccd1 hold5993/X sky130_fd_sc_hd__dlygate4sd3_1
X_12042_ _12267_/A _12042_/B vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 hold19/X vssd1 vssd1 vccd1 vccd1 input26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16850_ _18019_/CLK _16850_/D vssd1 vssd1 vccd1 vccd1 _16850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _17700_/CLK _15801_/D vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout770 fanout847/X vssd1 vssd1 vccd1 vccd1 fanout770/X sky130_fd_sc_hd__buf_4
XFILLER_0_137_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout781 _08147_/A vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__buf_4
X_16781_ _18014_/CLK _16781_/D vssd1 vssd1 vccd1 vccd1 _16781_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout792 fanout796/X vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__buf_2
XFILLER_0_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13993_ hold2804/X _13995_/A2 _13992_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _13993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15732_ _17703_/CLK _15732_/D vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ hold3280/X _12943_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18452_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _17207_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12875_ hold3149/X _12874_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__mux2_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _18452_/CLK _17402_/D vssd1 vssd1 vccd1 vccd1 _17402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _15169_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18382_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
X_11826_ _12213_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__or2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _17178_/CLK _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17523_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _17333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14545_ _15225_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14545_/X sky130_fd_sc_hd__or2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ hold4793/X _11667_/A _11756_/X vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10708_ hold5086/X _11198_/B _10707_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17264_ _17718_/CLK _17264_/D vssd1 vssd1 vccd1 vccd1 _17264_/Q sky130_fd_sc_hd__dfxtp_1
X_14476_ hold1823/X _14482_/A2 _14475_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14476_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11688_ _12234_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11688_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16215_ _17258_/CLK _16215_/D vssd1 vssd1 vccd1 vccd1 _16215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ hold1225/X _17596_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__mux2_1
X_10639_ _18461_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _16703_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17195_ _17195_/CLK _17195_/D vssd1 vssd1 vccd1 vccd1 _17195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _16148_/CLK _16146_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _15862_/Q _17573_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12309_ hold4645/X _12213_/A _12308_/X vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__a21oi_1
X_16077_ _16077_/CLK _16077_/D vssd1 vssd1 vccd1 vccd1 hold627/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _13289_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__and2_1
XFILLER_0_122_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3309 _12785_/X vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__dlygate4sd3_1
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2608 _07870_/X vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2619 _14209_/X vssd1 vssd1 vccd1 vccd1 _17905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07850_ hold2310/X _07865_/B _07849_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07850_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1907 _14915_/X vssd1 vssd1 vccd1 vccd1 _18242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1918 _08087_/X vssd1 vssd1 vccd1 vccd1 _15683_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1929 _15846_/Q vssd1 vssd1 vccd1 vccd1 hold1929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07781_ hold181/X vssd1 vssd1 vccd1 vccd1 _15219_/A sky130_fd_sc_hd__inv_8
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16979_ _17825_/CLK _16979_/D vssd1 vssd1 vccd1 vccd1 _16979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09520_ hold3835/X _10004_/B _09519_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18393_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09451_ _09456_/C _09456_/D _09450_/Y vssd1 vssd1 vccd1 vccd1 _16310_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_235_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08402_ hold2699/X _08440_/A2 _08401_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08402_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09382_ hold685/X _09392_/B _09362_/D hold429/X _09381_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08333_ _15557_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _15543_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08195_ _15529_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5201 _11260_/X vssd1 vssd1 vccd1 vccd1 _16910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5212 _17039_/Q vssd1 vssd1 vccd1 vccd1 hold5212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5223 _11452_/X vssd1 vssd1 vccd1 vccd1 _16974_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5234 _17254_/Q vssd1 vssd1 vccd1 vccd1 hold5234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5245 _10372_/X vssd1 vssd1 vccd1 vccd1 _16614_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4500 _13582_/X vssd1 vssd1 vccd1 vccd1 _17647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4511 _17675_/Q vssd1 vssd1 vccd1 vccd1 hold4511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5256 _16958_/Q vssd1 vssd1 vccd1 vccd1 hold5256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4522 _13465_/X vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5267 _11491_/X vssd1 vssd1 vccd1 vccd1 _16987_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4533 _17736_/Q vssd1 vssd1 vccd1 vccd1 hold4533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5278 _16978_/Q vssd1 vssd1 vccd1 vccd1 hold5278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5289 _09982_/X vssd1 vssd1 vccd1 vccd1 _16484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4544 _11866_/X vssd1 vssd1 vccd1 vccd1 _17112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4555 hold5873/X vssd1 vssd1 vccd1 vccd1 hold5874/A sky130_fd_sc_hd__buf_4
Xhold3810 _16799_/Q vssd1 vssd1 vccd1 vccd1 hold3810/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4566 _13771_/X vssd1 vssd1 vccd1 vccd1 _17710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3821 _17253_/Q vssd1 vssd1 vccd1 vccd1 hold3821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4577 hold5847/X vssd1 vssd1 vccd1 vccd1 hold5848/A sky130_fd_sc_hd__buf_4
XFILLER_0_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3832 _11233_/X vssd1 vssd1 vccd1 vccd1 _16901_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3843 _16367_/Q vssd1 vssd1 vccd1 vccd1 hold3843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4588 _15403_/X vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4599 _16524_/Q vssd1 vssd1 vccd1 vccd1 hold4599/X sky130_fd_sc_hd__buf_2
Xhold3854 _17722_/Q vssd1 vssd1 vccd1 vccd1 hold3854/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3865 _09937_/X vssd1 vssd1 vccd1 vccd1 _16469_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3876 _16468_/Q vssd1 vssd1 vccd1 vccd1 hold3876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3887 _09916_/X vssd1 vssd1 vccd1 vccd1 _16462_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_268_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18226_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3898 _16460_/Q vssd1 vssd1 vccd1 vccd1 hold3898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ hold2269/X _07978_/B _07978_/Y _08159_/A vssd1 vssd1 vccd1 vccd1 _07979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ hold3946/X _10004_/B _09717_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__o211a_1
X_10990_ hold4771/X _11177_/B _10989_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09649_ hold3900/X _10007_/B _09648_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09649_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _12738_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _17396_/D sky130_fd_sc_hd__and2_1
XFILLER_0_195_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ hold4431/X _12365_/B _11610_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11611_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ _12969_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _17373_/D sky130_fd_sc_hd__and2_1
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _14330_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ hold4311/X _11729_/B _11541_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14261_ hold1636/X _14272_/B _14260_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14261_/X
+ sky130_fd_sc_hd__o211a_1
X_11473_ hold5575/X _11768_/B _11472_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16000_ _18405_/CLK _16000_/D vssd1 vssd1 vccd1 vccd1 hold814/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13212_ hold4670/X _13211_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_2
X_10424_ hold2862/X _16632_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14192_ _15537_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14192_/X sky130_fd_sc_hd__or2_1
Xclkbuf_6_40_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_40_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13143_ _13199_/A1 _13141_/X _13142_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10355_ hold3122/X hold3874/X _10997_/S vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5790 output78/X vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_12
X_10286_ hold2520/X _16586_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__mux2_1
X_17951_ _18060_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _17560_/Q _17094_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ hold4205/X _13862_/B _12024_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12025_/X
+ sky130_fd_sc_hd__o211a_1
X_16902_ _17908_/CLK _16902_/D vssd1 vssd1 vccd1 vccd1 _16902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17882_ _17882_/CLK hold865/X vssd1 vssd1 vccd1 vccd1 hold864/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16833_ _18068_/CLK _16833_/D vssd1 vssd1 vccd1 vccd1 _16833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16764_ _17997_/CLK _16764_/D vssd1 vssd1 vccd1 vccd1 _16764_/Q sky130_fd_sc_hd__dfxtp_1
X_13976_ _15211_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15715_ _17746_/CLK _15715_/D vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfxtp_1
X_12927_ _12996_/A _12927_/B vssd1 vssd1 vccd1 vccd1 _17485_/D sky130_fd_sc_hd__and2_1
X_16695_ _18123_/CLK _16695_/D vssd1 vssd1 vccd1 vccd1 _16695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15646_ _17189_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_18434_ _18434_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _12921_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _17462_/D sky130_fd_sc_hd__and2_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18365_ _18397_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11809_ hold5134/X _13798_/A2 _11808_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15577_ _17245_/CLK _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12789_/A _12789_/B vssd1 vssd1 vccd1 vccd1 _17439_/D sky130_fd_sc_hd__and2_1
XFILLER_0_185_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17344_/CLK hold81/X vssd1 vssd1 vccd1 vccd1 _17316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ hold2886/X _14541_/B _14527_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14528_/X
+ sky130_fd_sc_hd__o211a_1
X_18296_ _18296_/CLK hold684/X vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17247_ _17903_/CLK _17247_/D vssd1 vssd1 vccd1 vccd1 _17247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14459_ _15193_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17178_ _17178_/CLK _17178_/D vssd1 vssd1 vccd1 vccd1 _17178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ _17313_/CLK _16129_/D vssd1 vssd1 vccd1 vccd1 hold647/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3106 _18276_/Q vssd1 vssd1 vccd1 vccd1 hold3106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3117 _14703_/X vssd1 vssd1 vccd1 vccd1 _18141_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08951_ hold174/X hold283/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3128 _17924_/Q vssd1 vssd1 vccd1 vccd1 hold3128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 _18349_/Q vssd1 vssd1 vccd1 vccd1 hold3139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2405 _18093_/Q vssd1 vssd1 vccd1 vccd1 hold2405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2416 _18365_/Q vssd1 vssd1 vccd1 vccd1 hold2416/X sky130_fd_sc_hd__dlygate4sd3_1
X_07902_ _15525_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07902_/X sky130_fd_sc_hd__or2_1
Xhold2427 _14035_/X vssd1 vssd1 vccd1 vccd1 _17821_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08882_ hold47/X hold409/X _08928_/S vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2438 _15705_/Q vssd1 vssd1 vccd1 vccd1 hold2438/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_361_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17113_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1704 _17805_/Q vssd1 vssd1 vccd1 vccd1 hold1704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _17965_/Q vssd1 vssd1 vccd1 vccd1 hold2449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1715 _09177_/X vssd1 vssd1 vccd1 vccd1 _16201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1726 _07813_/X vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ hold915/X _07881_/B vssd1 vssd1 vccd1 vccd1 _07833_/X sky130_fd_sc_hd__or2_1
Xhold1737 _15716_/Q vssd1 vssd1 vccd1 vccd1 hold1737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 becStatus[0] vssd1 vssd1 vccd1 vccd1 input1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1759 _17857_/Q vssd1 vssd1 vccd1 vccd1 hold1759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09503_ hold1389/X _13070_/A _10001_/C vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ hold819/X _16303_/Q vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09365_ _09386_/A _09365_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09369_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_93_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08316_ hold2727/X _08323_/B _08315_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ hold2206/X _09338_/A2 _09295_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_30 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_41 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_52 hold181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_63 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08247_ hold3017/X _08268_/B _08246_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08247_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_74 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 hold367/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 hold5854/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ hold1305/X _08209_/B _08177_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08178_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5020 _16832_/Q vssd1 vssd1 vccd1 vccd1 hold5020/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5031 _13717_/X vssd1 vssd1 vccd1 vccd1 _17692_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5042 _16787_/Q vssd1 vssd1 vccd1 vccd1 hold5042/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5053 _09538_/X vssd1 vssd1 vccd1 vccd1 _16336_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5064 _16558_/Q vssd1 vssd1 vccd1 vccd1 hold5064/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4330 _17717_/Q vssd1 vssd1 vccd1 vccd1 hold4330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_449_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5075 _11686_/X vssd1 vssd1 vccd1 vccd1 _17052_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ _10524_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__or2_1
Xhold4341 _11890_/X vssd1 vssd1 vccd1 vccd1 _17120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5086 _16758_/Q vssd1 vssd1 vccd1 vccd1 hold5086/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4352 _17702_/Q vssd1 vssd1 vccd1 vccd1 hold4352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5097 _12115_/X vssd1 vssd1 vccd1 vccd1 _17195_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4363 _11047_/X vssd1 vssd1 vccd1 vccd1 _16839_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4374 _17715_/Q vssd1 vssd1 vccd1 vccd1 hold4374/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4385 _16777_/Q vssd1 vssd1 vccd1 vccd1 hold4385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3640 _12375_/Y vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _13302_/A _10191_/A _10070_/X vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__a21oi_1
Xhold3651 _16644_/Q vssd1 vssd1 vccd1 vccd1 hold3651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4396 _13555_/X vssd1 vssd1 vccd1 vccd1 _17638_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3662 _16443_/Q vssd1 vssd1 vccd1 vccd1 hold3662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3673 _09751_/X vssd1 vssd1 vccd1 vccd1 _16407_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3684 _12378_/Y vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2950 _14749_/X vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3695 hold6025/X vssd1 vssd1 vccd1 vccd1 hold3695/X sky130_fd_sc_hd__clkbuf_2
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2961 _17789_/Q vssd1 vssd1 vccd1 vccd1 hold2961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2972 _14607_/X vssd1 vssd1 vccd1 vccd1 _18095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2983 _18278_/Q vssd1 vssd1 vccd1 vccd1 hold2983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2994 _09312_/X vssd1 vssd1 vccd1 vccd1 _16266_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13830_ hold5657/X _13734_/A _13829_/X vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13761_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10973_ _18016_/Q _16815_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15500_ _15500_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__and2_1
X_12712_ hold1203/X hold3410/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
X_16480_ _18202_/CLK _16480_/D vssd1 vssd1 vccd1 vccd1 _16480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13788_/A _13692_/B vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ hold830/X _15451_/A2 _09386_/D hold867/X _15426_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12643_ hold2959/X _17392_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18150_ _18208_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _15489_/A _15362_/B _15362_/C _15362_/D vssd1 vssd1 vccd1 vccd1 _15362_/X
+ sky130_fd_sc_hd__or4_1
X_12574_ hold1779/X hold3170/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17101_ _17199_/CLK _17101_/D vssd1 vssd1 vccd1 vccd1 _17101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ hold1534/X hold756/X _14312_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14313_/X
+ sky130_fd_sc_hd__o211a_1
X_18081_ _18113_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ hold2903/X hold4990/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15293_ _15490_/A1 _15285_/X _15292_/X _15490_/B1 _18403_/Q vssd1 vssd1 vccd1 vccd1
+ _15293_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17032_ _17129_/CLK _17032_/D vssd1 vssd1 vccd1 vccd1 _17032_/Q sky130_fd_sc_hd__dfxtp_1
X_14244_ _15193_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ hold2031/X _16976_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10407_ _11100_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14175_ hold2907/X _14198_/B _14174_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__o211a_1
X_11387_ hold2104/X hold4364/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _13126_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__or2_1
X_10338_ _10476_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13055_/C _13057_/B _17521_/Q vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__and3b_4
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17966_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_1
X_10269_ _11100_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12008_ hold982/X _17160_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_206_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17865_ _17897_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ _18017_/CLK _16816_/D vssd1 vssd1 vccd1 vccd1 _16816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17796_ _17935_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16747_ _18044_/CLK _16747_/D vssd1 vssd1 vccd1 vccd1 _16747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13959_ hold1454/X _13995_/A2 _13958_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16678_ _18078_/CLK _16678_/D vssd1 vssd1 vccd1 vccd1 _16678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18418_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15629_ _17257_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09150_ _15533_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__or2_1
X_18348_ _18380_/CLK hold748/X vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08101_ hold1477/X _08088_/B _08100_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _08101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18279_ _18377_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09081_ hold2304/X _09119_/A2 _09080_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08032_ hold2656/X _08033_/B _08031_/Y _08119_/A vssd1 vssd1 vccd1 vccd1 _08032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 input50/A vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_6
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_6
Xhold801 hold801/A vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold812 hold812/A vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 input70/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold834 hold834/A vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold845 hold845/A vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold856 hold856/A vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 hold878/A vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ hold1853/X hold3370/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__mux2_1
Xhold889 hold889/A vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2202 _07899_/X vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _08934_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _08963_/S sky130_fd_sc_hd__or2_2
XFILLER_0_200_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2213 _07864_/X vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2224 _08194_/X vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 _15108_/X vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 _18099_/Q vssd1 vssd1 vccd1 vccd1 hold2246/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1501 _17754_/Q vssd1 vssd1 vccd1 vccd1 hold1501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1512 _14315_/X vssd1 vssd1 vccd1 vccd1 _17955_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ _15454_/A hold709/X vssd1 vssd1 vccd1 vccd1 _16051_/D sky130_fd_sc_hd__and2_1
Xhold2257 _07981_/X vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2268 _08073_/X vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _15600_/Q vssd1 vssd1 vccd1 vccd1 hold1523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2279 _14149_/X vssd1 vssd1 vccd1 vccd1 _17876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _17954_/Q vssd1 vssd1 vccd1 vccd1 hold1534/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1545 _17884_/Q vssd1 vssd1 vccd1 vccd1 hold1545/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1556 _14785_/X vssd1 vssd1 vccd1 vccd1 _18181_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ _15515_/A _14972_/A hold999/A _14968_/A vssd1 vssd1 vccd1 vccd1 _07817_/D
+ sky130_fd_sc_hd__or4_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 _15729_/Q vssd1 vssd1 vccd1 vccd1 hold1567/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08796_ _08868_/B _08934_/A _13046_/D vssd1 vssd1 vccd1 vccd1 _08801_/S sky130_fd_sc_hd__or3_2
Xhold1578 _08300_/X vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 _17838_/Q vssd1 vssd1 vccd1 vccd1 hold1589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09417_ _07804_/A _09456_/A _15304_/A _09416_/X vssd1 vssd1 vccd1 vccd1 _09417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ hold246/A _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_0_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09279_ _15555_/A hold2752/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _12057_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11310_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ hold1670/X hold5234/X _13412_/S vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _11712_/A _11241_/B vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_283_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18053_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11172_ hold4660/X _11070_/A _11171_/X vssd1 vssd1 vccd1 vccd1 _11172_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_212_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18394_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4160 _17170_/Q vssd1 vssd1 vccd1 vccd1 hold4160/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ hold3712/X _10601_/B _10122_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10123_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4171 _17625_/Q vssd1 vssd1 vccd1 vccd1 hold4171/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4182 _09715_/X vssd1 vssd1 vccd1 vccd1 _16395_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _16087_/CLK _15980_/D vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__dfxtp_1
XTAP_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4193 _17124_/Q vssd1 vssd1 vccd1 vccd1 hold4193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3470 _17245_/Q vssd1 vssd1 vccd1 vccd1 hold3470/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14931_ hold1994/X _14946_/B _14930_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _14931_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10054_ _11194_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _16508_/D sky130_fd_sc_hd__nor2_1
Xhold3481 _12091_/X vssd1 vssd1 vccd1 vccd1 _17187_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3492 _17735_/Q vssd1 vssd1 vccd1 vccd1 hold3492/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2780 _15573_/Q vssd1 vssd1 vccd1 vccd1 hold2780/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _14862_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14862_/X sky130_fd_sc_hd__or2_1
X_17650_ _17650_/CLK _17650_/D vssd1 vssd1 vccd1 vccd1 _17650_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2791 _15738_/Q vssd1 vssd1 vccd1 vccd1 hold2791/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _18221_/CLK _16601_/D vssd1 vssd1 vccd1 vccd1 _16601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _13825_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _17724_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _17741_/CLK _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14793_ hold1344/X _14826_/B _14792_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14793_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16532_ _18152_/CLK _16532_/D vssd1 vssd1 vccd1 vccd1 _16532_/Q sky130_fd_sc_hd__dfxtp_1
X_13744_ _13838_/A _13856_/B _13743_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _17701_/D
+ sky130_fd_sc_hd__o211a_1
X_10956_ _11052_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16463_ _18342_/CLK _16463_/D vssd1 vssd1 vccd1 vccd1 _16463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ hold4525/X _13777_/A2 _13674_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13675_/X
+ sky130_fd_sc_hd__o211a_1
X_10887_ _11658_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15414_ _15414_/A _15414_/B vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__and2_1
X_18202_ _18202_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12626_ hold3323/X _12625_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__mux2_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _18395_/CLK _16394_/D vssd1 vssd1 vccd1 vccd1 _16394_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _18230_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
X_15345_ _15345_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12557_ hold3593/X _12556_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18064_ _18064_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_11508_ _12246_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11508_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15276_ _17331_/Q _15448_/B1 _15485_/B1 hold296/X vssd1 vssd1 vccd1 vccd1 _15276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12488_ _17337_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold180/X vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__buf_8
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17015_ _17902_/CLK _17015_/D vssd1 vssd1 vccd1 vccd1 _17015_/Q sky130_fd_sc_hd__dfxtp_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ hold1038/X _14216_/Y _14226_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _14227_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _11631_/A _11439_/B vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14158_ _15557_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _13108_/X hold4606/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14089_ hold2434/X _14094_/B _14088_/Y _15506_/A vssd1 vssd1 vccd1 vccd1 _14089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17917_ _18305_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08650_ _15324_/A hold644/X vssd1 vssd1 vccd1 vccd1 _15947_/D sky130_fd_sc_hd__and2_1
X_17848_ _17880_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08581_ _12408_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _15914_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_87_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16311_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17779_ _17875_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17478_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _15531_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ hold2848/X _09177_/A2 _09132_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09064_ _18459_/Q hold531/A vssd1 vssd1 vccd1 vccd1 hold532/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08015_ _15529_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 hold620/A vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 hold631/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold642 hold642/A vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold653 hold653/A vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold664 hold664/A vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 la_data_in[27] vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 hold697/A vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _10482_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__or2_1
Xhold2010 hold929/X vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _15604_/Q vssd1 vssd1 vccd1 vccd1 hold2021/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08917_ _12531_/A hold412/X vssd1 vssd1 vccd1 vccd1 _16076_/D sky130_fd_sc_hd__and2_1
Xhold2032 _14037_/X vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 _07949_/X vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09897_ _09918_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__or2_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2054 _18433_/Q vssd1 vssd1 vccd1 vccd1 hold2054/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _15880_/Q vssd1 vssd1 vccd1 vccd1 hold1320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2065 _17757_/Q vssd1 vssd1 vccd1 vccd1 hold2065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1331 hold6048/X vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__buf_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2076 _14484_/X vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _18289_/Q vssd1 vssd1 vccd1 vccd1 hold1342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2087 _18075_/Q vssd1 vssd1 vccd1 vccd1 hold2087/X sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ hold607/X hold901/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold902/A sky130_fd_sc_hd__mux2_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2098 _15832_/Q vssd1 vssd1 vccd1 vccd1 hold2098/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 _15712_/Q vssd1 vssd1 vccd1 vccd1 hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 _08077_/X vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _16223_/Q vssd1 vssd1 vccd1 vccd1 hold1375/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _09117_/X vssd1 vssd1 vccd1 vccd1 _16173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ hold578/X hold609/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1397 _17969_/Q vssd1 vssd1 vccd1 vccd1 hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ hold4823/X _11180_/B _10809_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10810_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ hold4998/X _11706_/A _11789_/X vssd1 vssd1 vccd1 vccd1 _11790_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ hold5633/X _11207_/B _10740_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ hold2295/X hold4269/X _13556_/S vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10672_ hold4238/X _11726_/B _10671_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _10672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12411_ hold346/X hold795/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold796/A sky130_fd_sc_hd__mux2_1
XFILLER_0_164_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13391_ hold2288/X hold3791/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_464_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15130_ hold1867/X _15165_/B _15129_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12342_ hold3724/X _12246_/A _12341_/X vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _15169_/A hold2273/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15062_/B sky130_fd_sc_hd__mux2_1
X_12273_ _12273_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14012_ _15519_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__or2_1
X_11224_ _12367_/A _11224_/B vssd1 vssd1 vccd1 vccd1 _16898_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _11158_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _16875_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ hold3236/X hold4687/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__mux2_1
XTAP_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_234_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15963_ _17314_/CLK _15963_/D vssd1 vssd1 vccd1 vccd1 hold482/A sky130_fd_sc_hd__dfxtp_1
X_11086_ hold4807/X _11180_/B _11085_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11086_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _17702_/CLK _17702_/D vssd1 vssd1 vccd1 vccd1 _17702_/Q sky130_fd_sc_hd__dfxtp_1
X_10037_ _16503_/Q _10037_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__and3_1
X_14914_ _15183_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14914_/X sky130_fd_sc_hd__or2_1
X_15894_ _17332_/CLK _15894_/D vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17728_/CLK _17633_/D vssd1 vssd1 vccd1 vccd1 _17633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14845_ hold1933/X _14880_/B _14844_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14776_ _15169_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14776_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17564_ _17724_/CLK _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_1
X_11988_ _13782_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16515_ _18266_/CLK _16515_/D vssd1 vssd1 vccd1 vccd1 _16515_/Q sky130_fd_sc_hd__dfxtp_1
X_13727_ hold1305/X _17696_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13728_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ hold5044/X _11216_/B _10938_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10939_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17495_ _17505_/CLK _17495_/D vssd1 vssd1 vccd1 vccd1 _17495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _18383_/CLK _16446_/D vssd1 vssd1 vccd1 vccd1 _16446_/Q sky130_fd_sc_hd__dfxtp_1
X_13658_ hold2199/X hold4315/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _13002_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _17379_/D sky130_fd_sc_hd__and2_1
X_16377_ _18350_/CLK _16377_/D vssd1 vssd1 vccd1 vccd1 _16377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13589_ hold1577/X _17650_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15328_ hold636/X _15484_/A2 _09392_/D hold320/X vssd1 vssd1 vccd1 vccd1 _15328_/X
+ sky130_fd_sc_hd__a22o_1
X_18116_ _18154_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_134_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17343_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5608 _10843_/X vssd1 vssd1 vccd1 vccd1 _16771_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5619 _16899_/Q vssd1 vssd1 vccd1 vccd1 hold5619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ hold537/X _15485_/A2 _15488_/A2 hold300/X _15258_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/C sky130_fd_sc_hd__a221o_1
X_18047_ _18337_/CLK _18047_/D vssd1 vssd1 vccd1 vccd1 _18047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4907 _16914_/Q vssd1 vssd1 vccd1 vccd1 hold4907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4918 _12016_/X vssd1 vssd1 vccd1 vccd1 _17162_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4929 _16734_/Q vssd1 vssd1 vccd1 vccd1 hold4929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ hold3986/X _10010_/B _09819_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09820_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout407 _14266_/B vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__buf_6
Xfanout418 _14052_/B vssd1 vssd1 vccd1 vccd1 _14042_/B sky130_fd_sc_hd__buf_6
XFILLER_0_22_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout429 _13054_/X vssd1 vssd1 vccd1 vccd1 _13309_/S sky130_fd_sc_hd__buf_12
XFILLER_0_201_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09751_ hold3672/X _10055_/B _09750_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08702_ _15344_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _15972_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09682_ hold4841/X _10571_/B _09681_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09682_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08633_ hold379/X hold562/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ hold256/X hold519/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08565_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ hold2599/X _08486_/B _08494_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09116_ _15557_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09047_ _12444_/A hold521/X vssd1 vssd1 vccd1 vccd1 _16140_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 hold450/A vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/A vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 hold483/A vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 hold494/A vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout930 _15211_/A vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__buf_12
Xfanout941 hold1019/X vssd1 vssd1 vccd1 vccd1 hold1020/A sky130_fd_sc_hd__buf_6
X_09949_ hold4833/X _10055_/B _09948_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09949_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_217_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _17496_/D sky130_fd_sc_hd__and2_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 hold1150/A vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 _18189_/Q vssd1 vssd1 vccd1 vccd1 hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ hold3774/X _12293_/B _11910_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _11911_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _15691_/Q vssd1 vssd1 vccd1 vccd1 hold1172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1183 _18074_/Q vssd1 vssd1 vccd1 vccd1 hold1183/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12975_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _17473_/D sky130_fd_sc_hd__and2_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _18321_/Q vssd1 vssd1 vccd1 vccd1 hold1194/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15131_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ hold5360/X _12031_/A2 _11841_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _11842_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14561_ hold915/X _14557_/Y _14560_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 hold916/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12340_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _17081_/D sky130_fd_sc_hd__nor2_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16320_/CLK _16300_/D vssd1 vssd1 vccd1 vccd1 _16300_/Q sky130_fd_sc_hd__dfxtp_1
X_13512_ _13800_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__or2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17280_/CLK _17280_/D vssd1 vssd1 vccd1 vccd1 _17280_/Q sky130_fd_sc_hd__dfxtp_1
X_10724_ hold2265/X hold3720/X _11204_/C vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__mux2_1
X_14492_ hold797/X _14487_/B _14491_/X _14360_/A vssd1 vssd1 vccd1 vccd1 hold798/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _17431_/CLK _16231_/D vssd1 vssd1 vccd1 vccd1 _16231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13443_ _13767_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10655_ hold1847/X _16709_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16162_ _17499_/CLK _16162_/D vssd1 vssd1 vccd1 vccd1 _16162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13374_ _13779_/A _13374_/B vssd1 vssd1 vccd1 vccd1 _13374_/X sky130_fd_sc_hd__or2_1
X_10586_ _16686_/Q _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__and3_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ _15221_/A _15113_/B vssd1 vssd1 vccd1 vccd1 _15113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12325_ _12340_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _17265_/D sky130_fd_sc_hd__nor2_1
X_16093_ _18399_/CLK _16093_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15044_ _15044_/A _15044_/B vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__and2_1
X_12256_ hold3978/X _12374_/B _12255_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12256_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_11207_ _16893_/Q _11207_/B _11768_/C vssd1 vssd1 vccd1 vccd1 _11207_/X sky130_fd_sc_hd__and3_1
X_12187_ hold4289/X _13877_/B _12186_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ _18071_/Q _16870_/Q _11150_/C vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16995_ _17870_/CLK _16995_/D vssd1 vssd1 vccd1 vccd1 _16995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15946_ _17293_/CLK _15946_/D vssd1 vssd1 vccd1 vccd1 hold636/A sky130_fd_sc_hd__dfxtp_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ hold1879/X hold3804/X _11168_/C vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _17745_/CLK _15877_/D vssd1 vssd1 vccd1 vccd1 _15877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _17739_/CLK _17616_/D vssd1 vssd1 vccd1 vccd1 _17616_/Q sky130_fd_sc_hd__dfxtp_1
X_14828_ _15221_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17547_ _18262_/CLK _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14759_ hold2465/X _14774_/B _14758_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_386_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17234_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08280_ _15559_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ _17478_/CLK _17478_/D vssd1 vssd1 vccd1 vccd1 _17478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_315_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18003_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16429_ _18380_/CLK _16429_/D vssd1 vssd1 vccd1 vccd1 _16429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5405 _17229_/Q vssd1 vssd1 vccd1 vccd1 hold5405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5416 _10681_/X vssd1 vssd1 vccd1 vccd1 _16717_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5427 _17244_/Q vssd1 vssd1 vccd1 vccd1 hold5427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5438 _11476_/X vssd1 vssd1 vccd1 vccd1 _16982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4704 _10987_/X vssd1 vssd1 vccd1 vccd1 _16819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5449 _16972_/Q vssd1 vssd1 vccd1 vccd1 hold5449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4715 _16883_/Q vssd1 vssd1 vccd1 vccd1 hold4715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4726 _10596_/Y vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4737 _16515_/Q vssd1 vssd1 vccd1 vccd1 hold4737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4748 _13863_/Y vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4759 _16374_/Q vssd1 vssd1 vccd1 vccd1 hold4759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _11584_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout215 _10019_/B vssd1 vssd1 vccd1 vccd1 _09832_/A2 sky130_fd_sc_hd__buf_4
Xfanout226 fanout246/X vssd1 vssd1 vccd1 vccd1 _10468_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout237 _10037_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_199_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09803_ hold2234/X _16425_/Q _10019_/C vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 _13623_/A vssd1 vssd1 vccd1 vccd1 _13800_/A sky130_fd_sc_hd__buf_4
XFILLER_0_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _14164_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__or2_1
Xfanout259 _11712_/A vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__buf_4
XFILLER_0_201_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09734_ hold844/X _16402_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_236_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ hold2654/X _16379_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ _12444_/A _08616_/B vssd1 vssd1 vccd1 vccd1 _15930_/D sky130_fd_sc_hd__and2_1
X_09596_ hold2981/X hold4024/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__mux2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _09063_/A hold619/X vssd1 vssd1 vccd1 vccd1 _15897_/D sky130_fd_sc_hd__and2_1
XFILLER_0_92_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08478_ _15211_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _10536_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_6_30_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_30_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_10371_ _10563_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ hold2015/X hold4917/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__mux2_1
Xhold5950 _17527_/Q vssd1 vssd1 vccd1 vccd1 hold5950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13090_ _17562_/Q _17096_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
Xhold5961 data_in[13] vssd1 vssd1 vccd1 vccd1 hold451/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5972 _16316_/Q vssd1 vssd1 vccd1 vccd1 hold5972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5983 _17514_/Q vssd1 vssd1 vccd1 vccd1 hold5983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5994 _18288_/Q vssd1 vssd1 vccd1 vccd1 hold5994/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12041_ hold2149/X hold4145/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__mux2_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 input26/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__buf_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout760 _13903_/A vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout771 _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__buf_4
X_15800_ _17667_/CLK _15800_/D vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout782 fanout796/X vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16780_ _18045_/CLK _16780_/D vssd1 vssd1 vccd1 vccd1 _16780_/Q sky130_fd_sc_hd__dfxtp_1
X_13992_ _15553_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout793 _14350_/A vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__buf_4
XFILLER_0_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12943_ hold2304/X hold3270/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__mux2_1
X_15731_ _17702_/CLK _15731_/D vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18450_ _18450_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _17113_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ hold975/X _17469_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17401_ _18438_/CLK _17401_/D vssd1 vssd1 vccd1 vccd1 _17401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ hold2447/X _14612_/B _14612_/Y _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14613_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11825_ hold1172/X hold4658/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__mux2_1
X_18381_ _18381_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
X_15593_ _17895_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17332_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 _17332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14544_ hold2349/X _14541_/B _14543_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14544_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _17076_/Q _11762_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _11756_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _11103_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _14529_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14475_/X sky130_fd_sc_hd__or2_1
X_17263_ _17263_/CLK _17263_/D vssd1 vssd1 vccd1 vccd1 _17263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ hold2160/X _17053_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13426_ hold4032/X _13802_/B _13425_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16214_ _17258_/CLK _16214_/D vssd1 vssd1 vccd1 vccd1 _16214_/Q sky130_fd_sc_hd__dfxtp_1
X_10638_ hold4649/X _10542_/A _10637_/X vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__a21oi_1
X_17194_ _17194_/CLK _17194_/D vssd1 vssd1 vccd1 vccd1 _17194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16145_ _17327_/CLK _16145_/D vssd1 vssd1 vccd1 vccd1 _16145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13357_ hold4547/X _13777_/A2 _13356_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _13357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10569_ hold4634/X _10563_/A _10568_/X vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _17260_/Q _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__and3_1
X_16076_ _17284_/CLK _16076_/D vssd1 vssd1 vccd1 vccd1 hold411/A sky130_fd_sc_hd__dfxtp_1
X_13288_ _13281_/X _13287_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_228_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15027_ _14116_/A hold2871/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__mux2_1
X_12239_ hold3021/X _17237_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2609 _15799_/Q vssd1 vssd1 vccd1 vccd1 hold2609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1908 _18183_/Q vssd1 vssd1 vccd1 vccd1 hold1908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1919 _16174_/Q vssd1 vssd1 vccd1 vccd1 hold1919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07780_ hold367/X vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_194_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16978_ _17884_/CLK _16978_/D vssd1 vssd1 vccd1 vccd1 _16978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15929_ _17347_/CLK _15929_/D vssd1 vssd1 vccd1 vccd1 hold613/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09450_ _09456_/C _09456_/D _09484_/B vssd1 vssd1 vccd1 vccd1 _09450_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_91_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08401_ _15515_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09381_ hold781/X _09386_/A _15479_/B1 hold701/X vssd1 vssd1 vccd1 vccd1 _09381_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08332_ hold2609/X _08323_/B _08331_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ hold2391/X _08263_/A2 _08262_/Y _08349_/A vssd1 vssd1 vccd1 vccd1 _08263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08194_ hold2223/X _08213_/B _08193_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _08194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5202 _16665_/Q vssd1 vssd1 vccd1 vccd1 hold5202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5213 _11551_/X vssd1 vssd1 vccd1 vccd1 _17007_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5224 _17064_/Q vssd1 vssd1 vccd1 vccd1 hold5224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5235 _12196_/X vssd1 vssd1 vccd1 vccd1 _17222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4501 _16432_/Q vssd1 vssd1 vccd1 vccd1 hold4501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5246 _17008_/Q vssd1 vssd1 vccd1 vccd1 hold5246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4512 _13570_/X vssd1 vssd1 vccd1 vccd1 _17643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5257 _11308_/X vssd1 vssd1 vccd1 vccd1 _16926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5268 _17590_/Q vssd1 vssd1 vccd1 vccd1 hold5268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4523 _16801_/Q vssd1 vssd1 vccd1 vccd1 hold4523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4534 _13753_/X vssd1 vssd1 vccd1 vccd1 _17704_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5279 _11368_/X vssd1 vssd1 vccd1 vccd1 _16946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4545 _17636_/Q vssd1 vssd1 vccd1 vccd1 hold4545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3800 _17398_/Q vssd1 vssd1 vccd1 vccd1 hold3800/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3811 _10831_/X vssd1 vssd1 vccd1 vccd1 _16767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4556 _15423_/X vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4567 _17708_/Q vssd1 vssd1 vccd1 vccd1 hold4567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3822 _12193_/X vssd1 vssd1 vccd1 vccd1 _17221_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4578 _15383_/X vssd1 vssd1 vccd1 vccd1 _15384_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3833 _16901_/Q vssd1 vssd1 vccd1 vccd1 hold3833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3844 _09535_/X vssd1 vssd1 vccd1 vccd1 _16335_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4589 hold5857/X vssd1 vssd1 vccd1 vccd1 hold5858/A sky130_fd_sc_hd__buf_6
Xhold3855 _13711_/X vssd1 vssd1 vccd1 vccd1 _17690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3866 _17661_/Q vssd1 vssd1 vccd1 vccd1 hold3866/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3877 _09838_/X vssd1 vssd1 vccd1 vccd1 _16436_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3888 _16500_/Q vssd1 vssd1 vccd1 vccd1 _10028_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3899 _09814_/X vssd1 vssd1 vccd1 vccd1 _16428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07978_ _15547_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07978_/Y sky130_fd_sc_hd__nand2_1
X_09717_ _09963_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__or2_1
XFILLER_0_198_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09648_ _09936_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__or2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_237_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18199_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10191_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09579_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11610_ _12246_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ hold3275/X _12589_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11541_ _11637_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14260_ _14529_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11694_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ _13210_/X _16919_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__mux2_1
X_10423_ hold3990/X _10631_/B _10422_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
X_14191_ hold1616/X _14202_/B _14190_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _14191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13142_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__or2_1
X_10354_ hold4002/X _10646_/B _10353_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5780 output73/X vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_12
X_13073_ _13073_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__and2_1
X_17950_ _18014_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5791 hold5934/X vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10285_ hold4162/X _10625_/B _10284_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10285_/X
+ sky130_fd_sc_hd__o211a_1
X_12024_ _12024_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__or2_1
X_16901_ _17907_/CLK _16901_/D vssd1 vssd1 vccd1 vccd1 _16901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17881_ _17975_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16832_ _18036_/CLK _16832_/D vssd1 vssd1 vccd1 vccd1 _16832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout590 _12751_/S vssd1 vssd1 vccd1 vccd1 _12772_/S sky130_fd_sc_hd__buf_6
XFILLER_0_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ _17996_/CLK _16763_/D vssd1 vssd1 vccd1 vccd1 _16763_/Q sky130_fd_sc_hd__dfxtp_1
X_13975_ hold1699/X _13995_/A2 _13974_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _13975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _17237_/CLK _15714_/D vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ hold3290/X _12925_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16694_ _18198_/CLK _16694_/D vssd1 vssd1 vccd1 vccd1 _16694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18433_ _18434_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _17157_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ hold3319/X _12856_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18364_/CLK hold904/X vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _13797_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15576_ _17244_/CLK _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ hold3317/X _12787_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/CLK _17315_/D vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14527_ _15099_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11739_ hold4697/X _11643_/A _11738_/X vssd1 vssd1 vccd1 vccd1 _11739_/Y sky130_fd_sc_hd__a21oi_1
X_18295_ _18327_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _17278_/CLK _17246_/D vssd1 vssd1 vccd1 vccd1 _17246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ hold2367/X _14482_/A2 _14457_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13409_ hold1744/X hold5268/X _13793_/S vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_226_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14389_ _15231_/A hold1701/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17177_ _17273_/CLK _17177_/D vssd1 vssd1 vccd1 vccd1 _17177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16128_ _16128_/CLK _16128_/D vssd1 vssd1 vccd1 vccd1 hold776/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3107 _14985_/X vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08950_ _12426_/A hold877/X vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__and2_1
XFILLER_0_228_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16059_ _18415_/CLK _16059_/D vssd1 vssd1 vccd1 vccd1 hold409/A sky130_fd_sc_hd__dfxtp_1
Xhold3118 _17997_/Q vssd1 vssd1 vccd1 vccd1 hold3118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3129 _14251_/X vssd1 vssd1 vccd1 vccd1 _17924_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07901_ hold1427/X _07918_/B _07900_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _07901_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2406 _14603_/X vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08881_ _15374_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _16058_/D sky130_fd_sc_hd__and2_1
Xhold2417 _15168_/X vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2428 _15680_/Q vssd1 vssd1 vccd1 vccd1 hold2428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2439 _15877_/Q vssd1 vssd1 vccd1 vccd1 hold2439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1705 _14003_/X vssd1 vssd1 vccd1 vccd1 _17805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 _17511_/Q vssd1 vssd1 vccd1 vccd1 hold1716/X sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ hold1585/X _07865_/B _07831_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07832_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1727 _09366_/A vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 _08154_/X vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 input1/X vssd1 vssd1 vccd1 vccd1 _13019_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ hold4024/X _10004_/B _09501_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09502_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_330_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09433_ _07804_/A _09477_/A _15344_/A hold825/X vssd1 vssd1 vccd1 vccd1 hold826/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09364_ _09366_/A _09364_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09364_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08315_ _15539_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09295_ _15517_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_31 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 hold181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _15525_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__or2_1
XANTENNA_64 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_75 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_86 hold367/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_97 hold5854/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08177_ hold915/X _08225_/B vssd1 vssd1 vccd1 vccd1 _08177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5010 _17195_/Q vssd1 vssd1 vccd1 vccd1 hold5010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5021 _10930_/X vssd1 vssd1 vccd1 vccd1 _16800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5032 _16450_/Q vssd1 vssd1 vccd1 vccd1 hold5032/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5043 _10795_/X vssd1 vssd1 vccd1 vccd1 _16755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5054 _16470_/Q vssd1 vssd1 vccd1 vccd1 hold5054/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5065 _10108_/X vssd1 vssd1 vccd1 vccd1 _16526_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4320 _11509_/X vssd1 vssd1 vccd1 vccd1 _16993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5076 _16438_/Q vssd1 vssd1 vccd1 vccd1 hold5076/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4331 _13696_/X vssd1 vssd1 vccd1 vccd1 _17685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5087 _10708_/X vssd1 vssd1 vccd1 vccd1 _16726_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4342 _17155_/Q vssd1 vssd1 vccd1 vccd1 hold4342/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5098 _16669_/Q vssd1 vssd1 vccd1 vccd1 hold5098/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4353 _13651_/X vssd1 vssd1 vccd1 vccd1 _17670_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4364 _16953_/Q vssd1 vssd1 vccd1 vccd1 hold4364/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3630 _13869_/Y vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4375 _13690_/X vssd1 vssd1 vccd1 vccd1 _17683_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10070_ _16514_/Q _10070_/B _10580_/C vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__and3_1
Xhold4386 _10765_/X vssd1 vssd1 vccd1 vccd1 _16745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3641 _17588_/Q vssd1 vssd1 vccd1 vccd1 hold3641/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4397 hold5863/X vssd1 vssd1 vccd1 vccd1 hold5864/A sky130_fd_sc_hd__buf_6
Xhold3652 _10366_/X vssd1 vssd1 vccd1 vccd1 _16612_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3663 _09763_/X vssd1 vssd1 vccd1 vccd1 _16411_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3674 _17429_/Q vssd1 vssd1 vccd1 vccd1 hold3674/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2940 _14027_/X vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3685 _16928_/Q vssd1 vssd1 vccd1 vccd1 hold3685/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2951 _18019_/Q vssd1 vssd1 vccd1 vccd1 hold2951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3696 _17414_/Q vssd1 vssd1 vccd1 vccd1 hold3696/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2962 _13969_/X vssd1 vssd1 vccd1 vccd1 _17789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 _18319_/Q vssd1 vssd1 vccd1 vccd1 hold2973/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_418_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17195_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_215_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2984 _14989_/X vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2995 _18280_/Q vssd1 vssd1 vccd1 vccd1 hold2995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13760_ hold2638/X hold4376/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10972_ hold5180/X _11159_/B _10971_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _12768_/A _12711_/B vssd1 vssd1 vccd1 vccd1 _17413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13691_ hold2674/X _17684_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13692_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15430_ hold712/X _09365_/B _09362_/D hold417/X _15428_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_167_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ _12759_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _17390_/D sky130_fd_sc_hd__and2_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _16300_/Q _15477_/A2 _15487_/B1 hold518/X _15360_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/D sky130_fd_sc_hd__a221o_1
X_12573_ _14362_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _17367_/D sky130_fd_sc_hd__and2_1
XFILLER_0_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17100_ _17260_/CLK _17100_/D vssd1 vssd1 vccd1 vccd1 _17100_/Q sky130_fd_sc_hd__dfxtp_1
X_11524_ hold5088/X _11617_/A2 _11523_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11524_/X
+ sky130_fd_sc_hd__o211a_1
X_14312_ _15207_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__or2_1
X_15292_ _15489_/A _15292_/B _15292_/C _15292_/D vssd1 vssd1 vccd1 vccd1 _15292_/X
+ sky130_fd_sc_hd__or4_1
X_18080_ _18112_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17031_ _18427_/CLK _17031_/D vssd1 vssd1 vccd1 vccd1 _17031_/Q sky130_fd_sc_hd__dfxtp_1
X_14243_ hold2113/X _14266_/B _14242_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ hold5314/X _12317_/B _11454_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ hold2865/X hold3668/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14174_ _15193_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ hold5587/X _11768_/B _11385_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11386_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _13124_/X hold4599/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__mux2_1
X_10337_ hold1962/X hold4803/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _17523_/Q _17522_/Q _13056_/C _13056_/D vssd1 vssd1 vccd1 vccd1 _13267_/S
+ sky130_fd_sc_hd__and4b_4
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _17997_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10268_ hold2850/X _16580_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10269_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ hold3837/X _12293_/B _12006_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _17896_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
X_10199_ hold3093/X _16557_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_159_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16815_ _18016_/CLK _16815_/D vssd1 vssd1 vccd1 vccd1 _16815_/Q sky130_fd_sc_hd__dfxtp_1
X_17795_ _18062_/CLK _17795_/D vssd1 vssd1 vccd1 vccd1 _17795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16746_ _18430_/CLK _16746_/D vssd1 vssd1 vccd1 vccd1 _16746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13958_ _15519_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ _12909_/A _12909_/B vssd1 vssd1 vccd1 vccd1 _17479_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16677_ _18233_/CLK _16677_/D vssd1 vssd1 vccd1 vccd1 _16677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ _07786_/Y _16286_/Q hold954/X _11057_/S vssd1 vssd1 vccd1 vccd1 _13889_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18416_ _18421_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15628_ _17444_/CLK _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18347_ _18379_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08100_ _14894_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _14910_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__or2_1
X_18278_ _18373_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ _15545_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput40 input40/A vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17229_ _17261_/CLK _17229_/D vssd1 vssd1 vccd1 vccd1 _17229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 input51/A vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xhold802 hold802/A vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold813 hold813/A vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold824 input70/X vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold835 hold835/A vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold857 hold857/A vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _13062_/A _10004_/B _09981_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09982_/X
+ sky130_fd_sc_hd__o211a_1
Xhold879 hold879/A vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ _15324_/A hold581/X vssd1 vssd1 vccd1 vccd1 _16084_/D sky130_fd_sc_hd__and2_1
Xhold2203 _17515_/Q vssd1 vssd1 vccd1 vccd1 hold2203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2214 _15770_/Q vssd1 vssd1 vccd1 vccd1 hold2214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2225 _15622_/Q vssd1 vssd1 vccd1 vccd1 hold2225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2236 _17835_/Q vssd1 vssd1 vccd1 vccd1 hold2236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2247 _14615_/X vssd1 vssd1 vccd1 vccd1 _18099_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ hold498/X hold708/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold709/A sky130_fd_sc_hd__mux2_1
XFILLER_0_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1502 _13896_/X vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _18126_/Q vssd1 vssd1 vccd1 vccd1 hold1513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2258 _17825_/Q vssd1 vssd1 vccd1 vccd1 hold2258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 _07913_/X vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 _15632_/Q vssd1 vssd1 vccd1 vccd1 hold2269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _14313_/X vssd1 vssd1 vccd1 vccd1 _17954_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07815_ _15523_/A _14910_/A _15519_/A _15517_/A vssd1 vssd1 vccd1 vccd1 _07817_/C
+ sky130_fd_sc_hd__or4_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1546 _14167_/X vssd1 vssd1 vccd1 vccd1 _17884_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ _13056_/C _13029_/A vssd1 vssd1 vccd1 vccd1 _13046_/D sky130_fd_sc_hd__nand2_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 _17872_/Q vssd1 vssd1 vccd1 vccd1 hold1557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1568 _08186_/X vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1579 _18199_/Q vssd1 vssd1 vccd1 vccd1 hold1579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09416_ _09438_/B _16294_/Q vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_220_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _09366_/A _09363_/B _09351_/B vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_191_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09278_ _12768_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _16250_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ hold203/X _15128_/A vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__or2_4
XFILLER_0_209_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ hold1949/X _16904_/Q _11711_/S vssd1 vssd1 vccd1 vccd1 _11241_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ _16881_/Q _11738_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__and3_1
XTAP_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4150 _13612_/X vssd1 vssd1 vccd1 vccd1 _17657_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10122_ _10488_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10122_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4161 _11944_/X vssd1 vssd1 vccd1 vccd1 _17138_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4172 _13420_/X vssd1 vssd1 vccd1 vccd1 _17593_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4183 hold5841/X vssd1 vssd1 vccd1 vccd1 hold5842/A sky130_fd_sc_hd__buf_4
XFILLER_0_235_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4194 _11806_/X vssd1 vssd1 vccd1 vccd1 _17092_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3460 _17205_/Q vssd1 vssd1 vccd1 vccd1 hold3460/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _15199_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14930_/X sky130_fd_sc_hd__or2_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10053_ _13254_/A _10467_/A _10052_/X vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__a21oi_1
Xhold3471 _12169_/X vssd1 vssd1 vccd1 vccd1 _17213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3482 _17649_/Q vssd1 vssd1 vccd1 vccd1 hold3482/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3493 _13750_/X vssd1 vssd1 vccd1 vccd1 _17703_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_252_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2770 _18192_/Q vssd1 vssd1 vccd1 vccd1 hold2770/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14861_ hold1977/X _14880_/B _14860_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14861_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2781 _07856_/X vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2792 _08204_/X vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _18220_/CLK _16600_/D vssd1 vssd1 vccd1 vccd1 _16600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13812_ hold4647/X _13716_/A _13811_/X vssd1 vssd1 vccd1 vccd1 _13812_/Y sky130_fd_sc_hd__a21oi_1
X_17580_ _17612_/CLK _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
X_14792_ _15131_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14792_/X sky130_fd_sc_hd__or2_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16531_ _18175_/CLK _16531_/D vssd1 vssd1 vccd1 vccd1 _16531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10955_ hold2570/X _16809_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__mux2_1
X_13743_ _13761_/A _13743_/B vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16462_ _18341_/CLK _16462_/D vssd1 vssd1 vccd1 vccd1 _16462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _13761_/A _13674_/B vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__or2_1
X_10886_ hold658/X hold5517/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18201_ _18201_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
X_15413_ _15490_/A1 _15405_/X _15412_/X _15490_/B1 hold5894/A vssd1 vssd1 vccd1 vccd1
+ _15413_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ hold2081/X _17386_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _18373_/CLK _16393_/D vssd1 vssd1 vccd1 vccd1 _16393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _18164_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ _15344_/A _15344_/B vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__and2_1
X_12556_ hold1547/X _17363_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ hold1975/X _16993_/Q _12365_/C vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18063_ _18063_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
X_12487_ hold56/X _12445_/A _12445_/B _12486_/X _12430_/A vssd1 vssd1 vccd1 vccd1
+ hold57/A sky130_fd_sc_hd__o311a_1
X_15275_ _15275_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _17892_/CLK _17014_/D vssd1 vssd1 vccd1 vccd1 _17014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14226_ hold926/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14226_/X sky130_fd_sc_hd__or2_1
X_11438_ hold2414/X hold4030/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14157_ hold2860/X _14148_/B _14156_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11369_ hold1873/X hold5537/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13108_ hold3262/X _13107_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__mux2_2
X_14088_ _15541_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_237_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ hold958/X _13039_/B vssd1 vssd1 vccd1 vccd1 hold959/A sky130_fd_sc_hd__and2_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17916_ _18014_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _17880_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ hold578/X hold648/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__mux2_1
X_17778_ _17907_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16729_ _17999_/CLK _16729_/D vssd1 vssd1 vccd1 vccd1 _16729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09201_ hold2527/X _09218_/B _09200_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _09201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09132_ _15515_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ _09063_/A hold187/X vssd1 vssd1 vccd1 vccd1 _16148_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ hold982/X _08029_/B _08013_/X _08353_/A vssd1 vssd1 vccd1 vccd1 hold983/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold610 hold610/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold621 hold716/X vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold643 hold643/A vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 hold654/A vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold665 hold665/A vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold676 hold676/A vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold687 hold687/A vssd1 vssd1 vccd1 vccd1 input56/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold698 hold698/A vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ hold887/X _16479_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__mux2_1
Xhold2000 _15767_/Q vssd1 vssd1 vccd1 vccd1 hold2000/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2011 input4/X vssd1 vssd1 vccd1 vccd1 hold930/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2022 _07921_/X vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08916_ hold263/X hold411/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold412/A sky130_fd_sc_hd__mux2_1
Xhold2033 _16271_/Q vssd1 vssd1 vccd1 vccd1 hold2033/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2044 _18460_/Q vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__buf_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _18367_/Q hold3351/X _10019_/C vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _09411_/X vssd1 vssd1 vccd1 vccd1 _16291_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2055 _15514_/X vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2066 _18011_/Q vssd1 vssd1 vccd1 vccd1 hold2066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _08506_/X vssd1 vssd1 vccd1 vccd1 _15880_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 _09409_/X vssd1 vssd1 vccd1 vccd1 _16290_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2077 _15756_/Q vssd1 vssd1 vccd1 vccd1 hold2077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _15011_/X vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2088 _14564_/X vssd1 vssd1 vccd1 vccd1 hold2088/X sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _12404_/A hold859/X vssd1 vssd1 vccd1 vccd1 _16042_/D sky130_fd_sc_hd__and2_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1354 hold1551/X vssd1 vssd1 vccd1 vccd1 hold1552/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2099 _08404_/X vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1365 _17949_/Q vssd1 vssd1 vccd1 vccd1 hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1376 _09223_/X vssd1 vssd1 vccd1 vccd1 _16223_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ _15482_/A hold267/X vssd1 vssd1 vccd1 vccd1 _16009_/D sky130_fd_sc_hd__and2_1
Xhold1387 _18373_/Q vssd1 vssd1 vccd1 vccd1 hold1387/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _18283_/Q vssd1 vssd1 vccd1 vccd1 hold1398/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ _11670_/A _10740_/B vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10671_ _11631_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _12412_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _17298_/D sky130_fd_sc_hd__and2_1
XFILLER_0_125_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13390_ hold4141/X _13868_/B _13389_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _13390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _17271_/Q _12365_/B _12365_/C vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ _15072_/A hold845/X vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12272_ hold2607/X _17248_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14011_ hold2153/X _14038_/B _14010_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14011_/X
+ sky130_fd_sc_hd__o211a_1
X_11223_ hold4919/X _11694_/A _11222_/X vssd1 vssd1 vccd1 vccd1 _11223_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_433_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17729_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ hold4903/X _11061_/A _11153_/X vssd1 vssd1 vccd1 vccd1 _11154_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ hold5344/X _10619_/B _10104_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10105_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _17315_/CLK _15962_/D vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__dfxtp_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _11100_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__or2_1
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ _17701_/CLK _17701_/D vssd1 vssd1 vccd1 vccd1 _17701_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3290 _17485_/Q vssd1 vssd1 vccd1 vccd1 hold3290/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ _11158_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _16502_/D sky130_fd_sc_hd__nor2_1
X_14913_ _14913_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14958_/B sky130_fd_sc_hd__or2_4
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15893_ _17339_/CLK _15893_/D vssd1 vssd1 vccd1 vccd1 hold494/A sky130_fd_sc_hd__dfxtp_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17632_ _17696_/CLK _17632_/D vssd1 vssd1 vccd1 vccd1 _17632_/Q sky130_fd_sc_hd__dfxtp_1
X_14844_ _15183_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17563_ _17723_/CLK _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775_ hold2524/X _14774_/B _14774_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11987_ hold1761/X _17153_/Q _13877_/C vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__mux2_1
X_16514_ _18265_/CLK _16514_/D vssd1 vssd1 vccd1 vccd1 _16514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13726_ hold5723/X _13829_/B _13725_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13726_/X
+ sky130_fd_sc_hd__o211a_1
X_10938_ _11121_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__or2_1
X_17494_ _17505_/CLK _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16445_ _18394_/CLK _16445_/D vssd1 vssd1 vccd1 vccd1 _16445_/Q sky130_fd_sc_hd__dfxtp_1
X_10869_ _11136_/A _10869_/B vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__or2_1
X_13657_ hold4393/X _13777_/A2 _13656_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _13657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ hold3577/X _12607_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _18287_/CLK _16376_/D vssd1 vssd1 vccd1 vccd1 _16376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ hold4505/X _13886_/B _13587_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13588_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ _18159_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15327_ _16141_/Q _15487_/A2 _15484_/B1 hold625/X _15326_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/B sky130_fd_sc_hd__a221o_1
X_12539_ hold3155/X _12538_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12539_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5609 _17079_/Q vssd1 vssd1 vccd1 vccd1 hold5609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18046_ _18046_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15258_ hold562/X _15484_/A2 _09392_/D hold407/X vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4908 _11751_/Y vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4919 _16738_/Q vssd1 vssd1 vccd1 vccd1 hold4919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ hold2618/X _14202_/B _14208_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14209_/X
+ sky130_fd_sc_hd__o211a_1
X_15189_ _15189_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_174_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18383_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout408 _14232_/Y vssd1 vssd1 vccd1 vccd1 _14266_/B sky130_fd_sc_hd__buf_8
Xfanout419 _14038_/B vssd1 vssd1 vccd1 vccd1 _14040_/B sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_103_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_238_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09750_ _09960_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08701_ hold568/X hold813/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__mux2_1
X_09681_ _10560_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08632_ _12416_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _15938_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08563_ _12424_/A hold439/X vssd1 vssd1 vccd1 vccd1 _15905_/D sky130_fd_sc_hd__and2_1
XFILLER_0_222_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08494_ _14726_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09115_ hold2553/X _09119_/A2 _09114_/X _12999_/A vssd1 vssd1 vccd1 vccd1 _09115_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_20_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_20_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ hold263/X hold520/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__mux2_1
XFILLER_0_241_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold440 hold440/A vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold451/A vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold473/A vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout920 hold972/X vssd1 vssd1 vccd1 vccd1 _14328_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout931 _15211_/A vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_217_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09948_ _09960_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__or2_1
Xfanout942 _15203_/A vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__buf_12
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _10191_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__or2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 la_data_in[22] vssd1 vssd1 vccd1 vccd1 hold1140/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 input37/X vssd1 vssd1 vccd1 vccd1 hold1151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _14803_/X vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _12288_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__or2_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1173 _18425_/Q vssd1 vssd1 vccd1 vccd1 hold1173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ hold3173/X _12889_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12890_/X sky130_fd_sc_hd__mux2_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _14562_/X vssd1 vssd1 vccd1 vccd1 hold1184/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _15078_/X vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _12024_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__or2_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14560_ hold690/X _14573_/B _18073_/Q vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__a21o_1
X_11772_ hold4905/X _12051_/A _11771_/X vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ hold5379/X _11201_/B _10722_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _10723_/X
+ sky130_fd_sc_hd__o211a_1
X_13511_ _15809_/Q _17624_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ hold559/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14491_/X sky130_fd_sc_hd__or2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16230_ _17431_/CLK _16230_/D vssd1 vssd1 vccd1 vccd1 _16230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ hold5463/X _11156_/B _10653_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10654_/X
+ sky130_fd_sc_hd__o211a_1
X_13442_ hold2867/X _17601_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16161_ _17499_/CLK _16161_/D vssd1 vssd1 vccd1 vccd1 _16161_/Q sky130_fd_sc_hd__dfxtp_1
X_13373_ hold1597/X _17578_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__mux2_1
X_10585_ _10603_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _16685_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15112_ hold885/X _15111_/B _15111_/Y _15066_/A vssd1 vssd1 vccd1 vccd1 hold886/A
+ sky130_fd_sc_hd__o211a_1
X_12324_ hold4871/X _12234_/A _12323_/X vssd1 vssd1 vccd1 vccd1 _12324_/Y sky130_fd_sc_hd__a21oi_1
X_16092_ _17304_/CLK _16092_/D vssd1 vssd1 vccd1 vccd1 hold876/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_1419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15043_ _15205_/A _18305_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ _13461_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12255_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ _12340_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _16892_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _13782_/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11137_ hold5493/X _11156_/B _11136_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _11137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16994_ _17862_/CLK _16994_/D vssd1 vssd1 vccd1 vccd1 _16994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15945_ _17327_/CLK _15945_/D vssd1 vssd1 vccd1 vccd1 hold405/A sky130_fd_sc_hd__dfxtp_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ hold5310/X _11201_/B _11067_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _11068_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ _16497_/Q _10019_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__and3_1
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _17737_/CLK _15876_/D vssd1 vssd1 vccd1 vccd1 _15876_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17647_/CLK _17615_/D vssd1 vssd1 vccd1 vccd1 _17615_/Q sky130_fd_sc_hd__dfxtp_1
X_14827_ hold2002/X _14826_/B _14826_/Y _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14827_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ _18294_/CLK _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14758_ _14758_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13709_ hold1515/X _17690_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17477_ _17478_/CLK _17477_/D vssd1 vssd1 vccd1 vccd1 _17477_/Q sky130_fd_sc_hd__dfxtp_1
X_14689_ hold3075/X _14720_/B _14688_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14689_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16428_ _18397_/CLK _16428_/D vssd1 vssd1 vccd1 vccd1 _16428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16359_ _18421_/CLK _16359_/D vssd1 vssd1 vccd1 vccd1 _16359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_355_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5406 _12121_/X vssd1 vssd1 vccd1 vccd1 _17197_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5417 _16989_/Q vssd1 vssd1 vccd1 vccd1 hold5417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5428 _12166_/X vssd1 vssd1 vccd1 vccd1 _17212_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5439 _16863_/Q vssd1 vssd1 vccd1 vccd1 hold5439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4705 _16409_/Q vssd1 vssd1 vccd1 vccd1 hold4705/X sky130_fd_sc_hd__dlygate4sd3_1
X_18029_ _18061_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4716 _11083_/X vssd1 vssd1 vccd1 vccd1 _16851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4727 _16594_/Q vssd1 vssd1 vccd1 vccd1 hold4727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4738 _09979_/X vssd1 vssd1 vccd1 vccd1 _16483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4749 _16477_/Q vssd1 vssd1 vccd1 vccd1 hold4749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout205 _11207_/B vssd1 vssd1 vccd1 vccd1 _11768_/B sky130_fd_sc_hd__clkbuf_8
Xfanout216 _10013_/B vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_238_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ hold3351/X _10013_/B _09801_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09802_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout227 _11095_/A2 vssd1 vssd1 vccd1 vccd1 _11198_/B sky130_fd_sc_hd__buf_4
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 _10037_/B vssd1 vssd1 vccd1 vccd1 _10577_/B sky130_fd_sc_hd__buf_2
XFILLER_0_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout249 _12288_/A vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__buf_4
X_07994_ hold203/X _14681_/A vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__or2_4
XFILLER_0_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09733_ hold4036/X _10010_/B _09732_/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 _09733_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ hold4843/X _10049_/B _09663_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09664_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ hold174/X hold546/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ hold4769/X _10601_/B _09594_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16320_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08546_ hold596/X hold618/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold619/A sky130_fd_sc_hd__mux2_1
XFILLER_0_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ hold1597/X _08486_/B _08476_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10370_ hold1931/X _16614_/Q _10580_/C vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09029_ _09055_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _16131_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5940 _17538_/Q vssd1 vssd1 vccd1 vccd1 hold5940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5951 _17526_/Q vssd1 vssd1 vccd1 vccd1 hold5951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5962 data_in[20] vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5973 data_in[18] vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ hold4217/X _13871_/B _12039_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _12040_/X
+ sky130_fd_sc_hd__o211a_1
Xhold270 input8/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5984 _18333_/Q vssd1 vssd1 vccd1 vccd1 hold5984/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5995 _15843_/Q vssd1 vssd1 vccd1 vccd1 hold5995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold292 hold20/X vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout750 fanout770/X vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout761 _13903_/A vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__buf_4
Xfanout772 _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13991_ hold1265/X _13986_/B _13990_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout783 _13941_/A vssd1 vssd1 vccd1 vccd1 _08127_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout794 _14350_/A vssd1 vssd1 vccd1 vccd1 _14548_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_217_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ _17732_/CLK _15730_/D vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12942_ _12996_/A _12942_/B vssd1 vssd1 vccd1 vccd1 _17490_/D sky130_fd_sc_hd__and2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _17269_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12912_/A _12873_/B vssd1 vssd1 vccd1 vccd1 _17467_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17400_ _18450_/CLK _17400_/D vssd1 vssd1 vccd1 vccd1 _17400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14612_ _14774_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__nand2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _18380_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11824_ hold4079/X _13811_/B _11823_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _11824_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _17210_/CLK _15592_/D vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17335_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _17331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _15169_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__or2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _12340_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _17075_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10706_ hold2496/X hold4632/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17262_ _17265_/CLK _17262_/D vssd1 vssd1 vccd1 vccd1 _17262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14474_ hold2917/X _14482_/A2 _14473_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ hold5074/X _12314_/B _11685_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11686_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16213_ _17258_/CLK _16213_/D vssd1 vssd1 vccd1 vccd1 _16213_/Q sky130_fd_sc_hd__dfxtp_1
X_13425_ _13713_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _13425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ _16703_/Q _10637_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17193_ _17257_/CLK _17193_/D vssd1 vssd1 vccd1 vccd1 _17193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _17330_/CLK _16144_/D vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10568_ _16680_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and3_1
X_13356_ _13776_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12307_ _12310_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _17259_/D sky130_fd_sc_hd__nor2_1
X_16075_ _17306_/CLK _16075_/D vssd1 vssd1 vccd1 vccd1 hold836/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ hold2443/X hold5393/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__mux2_1
X_13287_ _13311_/A1 _13285_/X _13286_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13287_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15026_ _15026_/A hold683/X vssd1 vssd1 vccd1 vccd1 hold684/A sky130_fd_sc_hd__and2_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12238_ hold4127/X _13868_/B _12237_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _12238_/X
+ sky130_fd_sc_hd__o211a_1
X_12169_ hold3470/X _13868_/B _12168_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12169_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1909 _14791_/X vssd1 vssd1 vccd1 vccd1 _18183_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16977_ _17855_/CLK _16977_/D vssd1 vssd1 vccd1 vccd1 _16977_/Q sky130_fd_sc_hd__dfxtp_1
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ _16148_/CLK _15928_/D vssd1 vssd1 vccd1 vccd1 hold371/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _17730_/CLK _15859_/D vssd1 vssd1 vccd1 vccd1 _15859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08400_ hold2715/X _08440_/A2 _08399_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08400_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09380_ hold722/X _09365_/B _09362_/A vssd1 vssd1 vccd1 vccd1 _09383_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_203_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ _15555_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08331_/X sky130_fd_sc_hd__or2_1
X_17529_ _17534_/CLK _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08262_ _14946_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08193_ _14862_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5203 _10429_/X vssd1 vssd1 vccd1 vccd1 _16633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5214 _17686_/Q vssd1 vssd1 vccd1 vccd1 hold5214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5225 _11626_/X vssd1 vssd1 vccd1 vccd1 _17032_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5236 _16632_/Q vssd1 vssd1 vccd1 vccd1 hold5236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4502 _09730_/X vssd1 vssd1 vccd1 vccd1 _16400_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5247 _11458_/X vssd1 vssd1 vccd1 vccd1 _16976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4513 _16828_/Q vssd1 vssd1 vccd1 vccd1 hold4513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5258 _17263_/Q vssd1 vssd1 vccd1 vccd1 hold5258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5269 _13315_/X vssd1 vssd1 vccd1 vccd1 _17558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4524 _10837_/X vssd1 vssd1 vccd1 vccd1 _16769_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4535 _16434_/Q vssd1 vssd1 vccd1 vccd1 hold4535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4546 _13453_/X vssd1 vssd1 vccd1 vccd1 _17604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3801 _17403_/Q vssd1 vssd1 vccd1 vccd1 hold3801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4557 _16898_/Q vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3812 _17127_/Q vssd1 vssd1 vccd1 vccd1 hold3812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3823 _16696_/Q vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4568 _13669_/X vssd1 vssd1 vccd1 vccd1 _17676_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4579 _17176_/Q vssd1 vssd1 vccd1 vccd1 hold4579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3834 _11713_/X vssd1 vssd1 vccd1 vccd1 _17061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3845 _17093_/Q vssd1 vssd1 vccd1 vccd1 hold3845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3856 _15995_/Q vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3867 _13528_/X vssd1 vssd1 vccd1 vccd1 _17629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3878 _16487_/Q vssd1 vssd1 vccd1 vccd1 hold3878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3889 _09934_/X vssd1 vssd1 vccd1 vccd1 _16468_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07977_ hold2504/X _07978_/B _07976_/Y _14149_/C1 vssd1 vssd1 vccd1 vccd1 _07977_/X
+ sky130_fd_sc_hd__o211a_1
X_09716_ hold1313/X _16396_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09717_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ hold1168/X _16373_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ hold1117/X _13270_/A _10190_/S vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ _15491_/A hold631/X vssd1 vssd1 vccd1 vccd1 _15889_/D sky130_fd_sc_hd__and2_1
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_277_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18078_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ hold2510/X hold4275/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_206_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18390_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ hold2573/X hold5561/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10422_ _10536_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__or2_1
X_13210_ _17577_/Q _17111_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _14529_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14190_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13141_ _13140_/X hold4687/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
X_10353_ _10998_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5770 output86/X vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_12
X_13072_ _13065_/X _13071_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17527_/D sky130_fd_sc_hd__o21a_1
Xhold5781 hold5921/X vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10284_ _10476_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5792 output76/X vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_12
X_12023_ hold2800/X _17165_/Q _12029_/S vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__mux2_1
X_16900_ _18426_/CLK _16900_/D vssd1 vssd1 vccd1 vccd1 _16900_/Q sky130_fd_sc_hd__dfxtp_1
X_17880_ _17880_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16831_ _18067_/CLK _16831_/D vssd1 vssd1 vccd1 vccd1 _16831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout580 _13057_/X vssd1 vssd1 vccd1 vccd1 _13306_/S sky130_fd_sc_hd__buf_8
Xfanout591 _12748_/S vssd1 vssd1 vccd1 vccd1 _12751_/S sky130_fd_sc_hd__buf_4
X_16762_ _17994_/CLK _16762_/D vssd1 vssd1 vccd1 vccd1 _16762_/Q sky130_fd_sc_hd__dfxtp_1
X_13974_ _14529_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15713_ _17585_/CLK _15713_/D vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12925_ _16149_/Q hold3264/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__mux2_1
X_16693_ _18219_/CLK _16693_/D vssd1 vssd1 vccd1 vccd1 _16693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ _18432_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
X_15644_ _17188_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ hold2848/X hold3314/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__mux2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18363_ _18363_/CLK hold963/X vssd1 vssd1 vccd1 vccd1 hold962/A sky130_fd_sc_hd__dfxtp_1
X_11807_ _15718_/Q hold3845/X _13412_/S vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15575_ _17590_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ hold2138/X _17440_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17314_ _17314_/CLK _17314_/D vssd1 vssd1 vccd1 vccd1 hold771/A sky130_fd_sc_hd__dfxtp_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ hold2542/X _14541_/B _14525_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14526_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18294_ _18294_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _17070_/Q _11738_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ _17245_/CLK _17245_/D vssd1 vssd1 vccd1 vccd1 _17245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _15191_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14457_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11669_ hold1626/X _17047_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ hold3474/X _13886_/B _13407_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17176_ _17872_/CLK _17176_/D vssd1 vssd1 vccd1 vccd1 _17176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ _14388_/A _14388_/B vssd1 vssd1 vccd1 vccd1 _17991_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _16127_/CLK _16127_/D vssd1 vssd1 vccd1 vccd1 _16127_/Q sky130_fd_sc_hd__dfxtp_1
X_13339_ hold5138/X _13817_/B _13338_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ _16081_/CLK _16058_/D vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__dfxtp_1
Xhold3108 _16157_/Q vssd1 vssd1 vccd1 vccd1 hold3108/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3119 _14402_/X vssd1 vssd1 vccd1 vccd1 _17997_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ hold5994/X _15004_/B hold980/X _15070_/A vssd1 vssd1 vccd1 vccd1 hold981/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07900_ _14517_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07900_/X sky130_fd_sc_hd__or2_1
Xhold2407 _18121_/Q vssd1 vssd1 vccd1 vccd1 hold2407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08880_ hold17/X hold339/X _08928_/S vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__mux2_1
Xhold2418 _16274_/Q vssd1 vssd1 vccd1 vccd1 hold2418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2429 _08081_/X vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1706 _15755_/Q vssd1 vssd1 vccd1 vccd1 hold1706/X sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ _15509_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07831_/X sky130_fd_sc_hd__or2_1
Xhold1717 _13006_/X vssd1 vssd1 vccd1 vccd1 _17511_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1728 _09401_/X vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _18233_/Q vssd1 vssd1 vccd1 vccd1 hold1739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09501_ _09987_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ hold819/X _16302_/Q vssd1 vssd1 vccd1 vccd1 hold825/A sky130_fd_sc_hd__or2_1
XFILLER_0_172_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _09366_/A _09363_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09363_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_370_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17707_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08314_ hold2896/X _08323_/B _08313_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08314_/X
+ sky130_fd_sc_hd__o211a_1
X_09294_ hold2901/X _09338_/A2 _09293_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_10 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_32 _17524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08245_ hold1662/X _08263_/A2 _08244_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_43 _15513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 hold181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_65 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 hold367/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ hold1164/X _08209_/B _08175_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5000 _16637_/Q vssd1 vssd1 vccd1 vccd1 hold5000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5011 _12019_/X vssd1 vssd1 vccd1 vccd1 _17163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5022 _17259_/Q vssd1 vssd1 vccd1 vccd1 hold5022/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5033 _09784_/X vssd1 vssd1 vccd1 vccd1 _16418_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5044 _16835_/Q vssd1 vssd1 vccd1 vccd1 hold5044/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5055 _09844_/X vssd1 vssd1 vccd1 vccd1 _16438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4310 _13648_/X vssd1 vssd1 vccd1 vccd1 _17669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5066 _16845_/Q vssd1 vssd1 vccd1 vccd1 hold5066/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4321 _17637_/Q vssd1 vssd1 vccd1 vccd1 hold4321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4332 _16993_/Q vssd1 vssd1 vccd1 vccd1 hold4332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5077 _09748_/X vssd1 vssd1 vccd1 vccd1 _16406_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4343 _11899_/X vssd1 vssd1 vccd1 vccd1 _17123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5088 _17030_/Q vssd1 vssd1 vccd1 vccd1 hold5088/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5099 _10441_/X vssd1 vssd1 vccd1 vccd1 _16637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4354 _16959_/Q vssd1 vssd1 vccd1 vccd1 hold4354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3620 _09559_/X vssd1 vssd1 vccd1 vccd1 _16343_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4365 _11293_/X vssd1 vssd1 vccd1 vccd1 _16921_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3631 _16377_/Q vssd1 vssd1 vccd1 vccd1 hold3631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4376 _17707_/Q vssd1 vssd1 vccd1 vccd1 hold4376/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4387 _16808_/Q vssd1 vssd1 vccd1 vccd1 hold4387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3642 _13884_/Y vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3653 _16379_/Q vssd1 vssd1 vccd1 vccd1 hold3653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4398 _09385_/X vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3664 _16888_/Q vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3675 _12758_/X vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2930 _07911_/X vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2941 _18108_/Q vssd1 vssd1 vccd1 vccd1 hold2941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3686 _11793_/Y vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2952 _14446_/X vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3697 _17577_/Q vssd1 vssd1 vccd1 vccd1 hold3697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 _18332_/Q vssd1 vssd1 vccd1 vccd1 hold2963/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2974 _17928_/Q vssd1 vssd1 vccd1 vccd1 hold2974/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2985 _17843_/Q vssd1 vssd1 vccd1 vccd1 hold2985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2996 _14993_/X vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _11064_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10971_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_458_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17420_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12710_ hold3781/X _12709_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13690_ hold4374/X _13880_/B _13689_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12641_ hold4157/X _12640_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ hold582/X _15486_/A2 _09357_/B hold396/X vssd1 vssd1 vccd1 vccd1 _15360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ hold3498/X _12571_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ hold1281/X hold756/X _14310_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _14311_/X
+ sky130_fd_sc_hd__o211a_1
X_11523_ _11712_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__or2_1
X_15291_ _16293_/Q _15477_/A2 _15487_/B1 hold356/X _15290_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _17876_/CLK _17030_/D vssd1 vssd1 vccd1 vccd1 _17030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _14403_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ _12285_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10405_ hold5393/X _10619_/B _10404_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14173_ hold2132/X _14198_/B _14172_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14173_/X
+ sky130_fd_sc_hd__o211a_1
X_11385_ _11694_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13124_ hold4911/X _13123_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10336_ hold4839/X _10649_/B _10335_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _17523_/Q _13056_/C _13055_/C _17522_/Q vssd1 vssd1 vccd1 vccd1 _13055_/X
+ sky130_fd_sc_hd__or4b_4
X_10267_ hold4805/X _10649_/B _10266_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17932_ _18050_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _12288_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__or2_1
X_17863_ _17863_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ hold4741/X _10598_/B _10197_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16814_ _18016_/CLK _16814_/D vssd1 vssd1 vccd1 vccd1 _16814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17794_ _17892_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16745_ _18012_/CLK _16745_/D vssd1 vssd1 vccd1 vccd1 _16745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13957_ hold2337/X _13995_/A2 _13956_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _13957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_199_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12908_ hold3391/X _12907_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12909_/B sky130_fd_sc_hd__mux2_1
X_16676_ _18232_/CLK _16676_/D vssd1 vssd1 vccd1 vccd1 _16676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _17749_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_159_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17320_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18415_ _18415_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_15627_ _17194_/CLK _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ hold3407/X _12838_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12840_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18346_ _18346_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15558_ hold1807/X _15560_/A2 _15557_/X _12654_/A vssd1 vssd1 vccd1 vccd1 _15558_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ _14974_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__or2_1
X_18277_ _18381_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15489_ _15489_/A _15489_/B _15489_/C _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_115_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ hold2017/X _08029_/B _08029_/Y _08161_/A vssd1 vssd1 vccd1 vccd1 _08030_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ _17260_/CLK _17228_/D vssd1 vssd1 vccd1 vccd1 _17228_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 input30/A vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput41 input41/A vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold814 hold814/A vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ _17194_/CLK _17159_/D vssd1 vssd1 vccd1 vccd1 _17159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold825 hold825/A vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold836 hold836/A vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold847 hold847/A vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 hold869/A vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _09987_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08932_ hold150/X hold580/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold581/A sky130_fd_sc_hd__mux2_1
XFILLER_0_209_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2204 _13014_/X vssd1 vssd1 vccd1 vccd1 _17515_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 _08271_/X vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_239_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2226 _07959_/X vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2237 _14065_/X vssd1 vssd1 vccd1 vccd1 _17835_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ _12418_/A hold800/X vssd1 vssd1 vccd1 vccd1 _16050_/D sky130_fd_sc_hd__and2_1
Xhold1503 _17940_/Q vssd1 vssd1 vccd1 vccd1 hold1503/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2248 _15567_/Q vssd1 vssd1 vccd1 vccd1 hold2248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 _14671_/X vssd1 vssd1 vccd1 vccd1 _18126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2259 _14043_/X vssd1 vssd1 vccd1 vccd1 _17825_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1525 _17778_/Q vssd1 vssd1 vccd1 vccd1 hold1525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07814_ _15105_/A _15103_/A _15535_/A _15099_/A vssd1 vssd1 vccd1 vccd1 _07817_/B
+ sky130_fd_sc_hd__or4_1
Xhold1536 _15827_/Q vssd1 vssd1 vccd1 vccd1 hold1536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _16261_/Q vssd1 vssd1 vccd1 vccd1 hold1547/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08794_ _15482_/A hold177/X vssd1 vssd1 vccd1 vccd1 _16017_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1558 _14141_/X vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1569 _18152_/Q vssd1 vssd1 vccd1 vccd1 hold1569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _07804_/A _09456_/B _15264_/A _09414_/X vssd1 vssd1 vccd1 vccd1 _09415_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09346_ hold367/A hold181/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__or3_2
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _15553_/A hold2784/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ hold203/X _15128_/A vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11170_ _12310_/A _11170_/B vssd1 vssd1 vccd1 vccd1 _16880_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4140 _12689_/X vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10121_ hold2280/X _16531_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4151 _17250_/Q vssd1 vssd1 vccd1 vccd1 hold4151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4162 _16617_/Q vssd1 vssd1 vccd1 vccd1 hold4162/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4173 _17150_/Q vssd1 vssd1 vccd1 vccd1 hold4173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4184 _15273_/X vssd1 vssd1 vccd1 vccd1 _15274_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4195 _16678_/Q vssd1 vssd1 vccd1 vccd1 hold4195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3450 _17213_/Q vssd1 vssd1 vccd1 vccd1 hold3450/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ _10052_/A _10070_/B _10190_/S vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__and3_1
Xhold3461 _12049_/X vssd1 vssd1 vccd1 vccd1 _17173_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3472 _17365_/Q vssd1 vssd1 vccd1 vccd1 hold3472/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3483 _13492_/X vssd1 vssd1 vccd1 vccd1 _17617_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3494 _17184_/Q vssd1 vssd1 vccd1 vccd1 hold3494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2760 _14279_/X vssd1 vssd1 vccd1 vccd1 _17938_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14860_ _15199_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__or2_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2771 _14809_/X vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2782 _18443_/Q vssd1 vssd1 vccd1 vccd1 hold2782/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2793 _15595_/Q vssd1 vssd1 vccd1 vccd1 hold2793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _17724_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _13811_/X sky130_fd_sc_hd__and3_1
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ hold1908/X _14826_/B _14790_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14791_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_292_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17825_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _18234_/CLK _16530_/D vssd1 vssd1 vccd1 vccd1 _16530_/Q sky130_fd_sc_hd__dfxtp_1
X_13742_ hold2333/X hold4309/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13743_/B sky130_fd_sc_hd__mux2_1
X_10954_ hold4346/X _11147_/B _10953_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_221_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18209_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16461_ _18276_/CLK _16461_/D vssd1 vssd1 vccd1 vccd1 _16461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13673_ hold2375/X _17678_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13674_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ hold3926/X _11738_/B _10884_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10885_/X
+ sky130_fd_sc_hd__o211a_1
X_18200_ _18200_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15412_ _15489_/A _15412_/B _15412_/C _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ _12780_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _17384_/D sky130_fd_sc_hd__and2_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _18303_/CLK _16392_/D vssd1 vssd1 vccd1 vccd1 _16392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18131_ _18131_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15343_ _15490_/A1 _15335_/X _15342_/X _15490_/B1 hold5836/A vssd1 vssd1 vccd1 vccd1
+ _15343_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _13002_/A _12555_/B vssd1 vssd1 vccd1 vccd1 _17361_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ hold4293/X _11801_/B _11505_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__o211a_1
X_18062_ _18062_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
X_15274_ _15344_/A _15274_/B vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__and2_1
XFILLER_0_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _17336_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17013_ _17901_/CLK _17013_/D vssd1 vssd1 vccd1 vccd1 _17013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14225_ hold1869/X _14216_/Y _14224_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _14225_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ hold3912/X _11726_/B _11436_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _15229_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11368_ hold5278/X _11738_/B _11367_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11368_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _13106_/X hold5911/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
X_10319_ hold2826/X _16597_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14087_ hold2725/X _14094_/B _14086_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _14087_/X
+ sky130_fd_sc_hd__o211a_1
X_11299_ hold5320/X _11747_/B _11298_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13038_ _13048_/A _13034_/X _17523_/Q vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__a21o_1
X_17915_ _18429_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _18427_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_309_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17966_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_234_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ hold2983/X hold514/X _14988_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _14989_/X
+ sky130_fd_sc_hd__o211a_1
X_17777_ _17777_/CLK _17777_/D vssd1 vssd1 vccd1 vccd1 _17777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ _18026_/CLK _16728_/D vssd1 vssd1 vccd1 vccd1 _16728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _18215_/CLK _16659_/D vssd1 vssd1 vccd1 vccd1 _16659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09200_ _15529_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09131_ hold2757/X _09177_/A2 _09130_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09131_/X
+ sky130_fd_sc_hd__o211a_1
X_18329_ _18391_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_6_10_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_10_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ hold150/X hold186/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_96_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08013_ hold944/X _08045_/B vssd1 vssd1 vccd1 vccd1 _08013_/X sky130_fd_sc_hd__or2_1
Xhold600 hold805/X vssd1 vssd1 vccd1 vccd1 hold806/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 hold611/A vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17507_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold622 hold718/X vssd1 vssd1 vccd1 vccd1 hold719/A sky130_fd_sc_hd__buf_6
Xhold633 hold633/A vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold644 hold644/A vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold655 hold655/A vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold666 hold666/A vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold677 hold677/A vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold688 input56/X vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__buf_1
Xhold699 hold699/A vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _10058_/A _10034_/B _09963_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09964_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2001 _08265_/X vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2012 _07811_/X vssd1 vssd1 vccd1 vccd1 hold2012/X sky130_fd_sc_hd__buf_1
XFILLER_0_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08915_ _12426_/A hold837/X vssd1 vssd1 vccd1 vccd1 _16075_/D sky130_fd_sc_hd__and2_1
Xhold2023 _17874_/Q vssd1 vssd1 vccd1 vccd1 hold2023/X sky130_fd_sc_hd__dlygate4sd3_1
X_09895_ hold3878/X _10013_/B _09894_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09895_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2034 _09322_/X vssd1 vssd1 vccd1 vccd1 _16271_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _07807_/X vssd1 vssd1 vccd1 vccd1 hold2045/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 hold1400/X vssd1 vssd1 vccd1 vccd1 hold1401/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 _15884_/Q vssd1 vssd1 vccd1 vccd1 hold2056/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _16249_/Q vssd1 vssd1 vccd1 vccd1 hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 _15715_/Q vssd1 vssd1 vccd1 vccd1 hold1322/X sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ hold228/X hold858/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold859/A sky130_fd_sc_hd__mux2_1
Xhold2067 _14430_/X vssd1 vssd1 vccd1 vccd1 _18011_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1333 hold1438/X vssd1 vssd1 vccd1 vccd1 hold1439/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 _08243_/X vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 _18184_/Q vssd1 vssd1 vccd1 vccd1 hold1344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2089 _14565_/X vssd1 vssd1 vccd1 vccd1 _18075_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1355 hold1553/X vssd1 vssd1 vccd1 vccd1 hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _14303_/X vssd1 vssd1 vccd1 vccd1 _17949_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1377 _17844_/Q vssd1 vssd1 vccd1 vccd1 hold1377/X sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ hold263/X hold266/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1388 _15186_/X vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _14999_/X vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ hold2453/X hold3262/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09329_ _15551_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _12340_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _17270_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _12365_/A _12365_/B _12270_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _12271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14010_ _14403_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__or2_1
X_11222_ _11222_/A _11768_/B _11768_/C vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__and3_1
XFILLER_0_222_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _11153_/A _11156_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ _10524_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__or2_1
XTAP_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15961_ _16128_/CLK _15961_/D vssd1 vssd1 vccd1 vccd1 hold881/A sky130_fd_sc_hd__dfxtp_1
X_11084_ hold1450/X hold4771/X _11192_/C vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__mux2_1
XTAP_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3280 _17491_/Q vssd1 vssd1 vccd1 vccd1 hold3280/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _13206_/A _09963_/A _10034_/X vssd1 vssd1 vccd1 vccd1 _10035_/Y sky130_fd_sc_hd__a21oi_1
X_14912_ _14913_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__nor2_2
X_17700_ _17700_/CLK _17700_/D vssd1 vssd1 vccd1 vccd1 _17700_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3291 _12926_/X vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15892_ _16148_/CLK _15892_/D vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__dfxtp_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2590 _15610_/Q vssd1 vssd1 vccd1 vccd1 hold2590/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_402_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ _14843_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14892_/B sky130_fd_sc_hd__or2_4
X_17631_ _17730_/CLK _17631_/D vssd1 vssd1 vccd1 vccd1 _17631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ _17722_/CLK _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_1
X_14774_ _14774_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11986_ hold3494/X _12274_/A2 _11985_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11986_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16513_ _16517_/CLK _16513_/D vssd1 vssd1 vccd1 vccd1 _16513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13725_ _13734_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ hold3080/X _16803_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__mux2_1
X_17493_ _17509_/CLK _17493_/D vssd1 vssd1 vccd1 vccd1 _17493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16444_ _18379_/CLK _16444_/D vssd1 vssd1 vccd1 vccd1 _16444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13746_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__or2_1
X_10868_ hold1903/X hold5336/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ hold1877/X _17380_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16375_ _18390_/CLK _16375_/D vssd1 vssd1 vccd1 vccd1 _16375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13587_ _13779_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__or2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ hold2583/X hold5130/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__mux2_1
X_18114_ _18224_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15326_ _17336_/Q _15448_/B1 _15485_/B1 hold169/X vssd1 vssd1 vccd1 vccd1 _15326_/X
+ sky130_fd_sc_hd__a22o_1
X_12538_ hold1327/X _17357_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18045_ _18045_/CLK hold871/X vssd1 vssd1 vccd1 vccd1 hold870/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15257_ hold616/X _15487_/A2 _15484_/B1 hold284/X _15256_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/B sky130_fd_sc_hd__a221o_1
X_12469_ hold361/X _12445_/A _12445_/B _12468_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold24/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4909 _16596_/Q vssd1 vssd1 vccd1 vccd1 hold4909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14208_ _14726_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15188_ hold856/X _15219_/B _15187_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 hold857/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ hold1763/X _14142_/B _14138_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout409 _14206_/B vssd1 vssd1 vccd1 vccd1 _14214_/B sky130_fd_sc_hd__buf_8
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ _15304_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _15971_/D sky130_fd_sc_hd__and2_1
XFILLER_0_59_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09680_ hold1072/X hold4731/X _10571_/C vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_143_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08631_ hold256/X hold410/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08632_/B sky130_fd_sc_hd__mux2_1
X_17829_ _17891_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08562_ hold346/X hold438/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__mux2_1
XFILLER_0_234_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08493_ hold1538/X _08486_/B _08492_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _08493_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09114_ _15555_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09045_ _15364_/A hold638/X vssd1 vssd1 vccd1 vccd1 _16139_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold441 hold441/A vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold452 hold73/X vssd1 vssd1 vccd1 vccd1 input9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold485 hold522/X vssd1 vssd1 vccd1 vccd1 hold523/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold496 hold76/X vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout910 _15121_/A vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__buf_12
XFILLER_0_239_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout921 hold972/X vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__buf_12
X_09947_ hold1452/X hold3345/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__mux2_1
Xfanout932 hold1355/X vssd1 vssd1 vccd1 vccd1 hold1356/A sky130_fd_sc_hd__buf_6
XFILLER_0_216_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout943 _15203_/A vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09878_ hold1573/X hold5032/X _10580_/C vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__mux2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _15731_/Q vssd1 vssd1 vccd1 vccd1 hold1130/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 hold1141/A vssd1 vssd1 vccd1 vccd1 input51/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _12436_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _16033_/D sky130_fd_sc_hd__and2_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 hold1152/A vssd1 vssd1 vccd1 vccd1 hold1152/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1163 _15717_/Q vssd1 vssd1 vccd1 vccd1 hold1163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1174 _18225_/Q vssd1 vssd1 vccd1 vccd1 hold1174/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _14563_/X vssd1 vssd1 vccd1 vccd1 _18074_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1196 _16241_/Q vssd1 vssd1 vccd1 vccd1 hold1196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ hold1040/X hold4719/X _13793_/S vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _17081_/Q _12338_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__and3_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13510_ hold3938/X _13802_/B _13509_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ _11106_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ hold2581/X _14487_/B _14489_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _14490_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ hold5761/X _13832_/B _13440_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13441_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _11136_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16160_ _17496_/CLK _16160_/D vssd1 vssd1 vccd1 vccd1 _16160_/Q sky130_fd_sc_hd__dfxtp_1
X_13372_ hold4356/X _13880_/B _13371_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ hold4627/X _10488_/A _10583_/X vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15111_ _15219_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _17265_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and3_1
X_16091_ _17299_/CLK _16091_/D vssd1 vssd1 vccd1 vccd1 hold846/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15042_ _15473_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ hold1367/X _17242_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ hold3720/X _11658_/A _11204_/X vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12185_ hold2399/X hold3480/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11136_ _11136_/A _11136_/B vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__or2_1
X_16993_ _17871_/CLK _16993_/D vssd1 vssd1 vccd1 vccd1 _16993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ _17299_/CLK _15944_/D vssd1 vssd1 vccd1 vccd1 hold838/A sky130_fd_sc_hd__dfxtp_1
X_11067_ _11106_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__or2_1
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _11158_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _16496_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_222_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15875_ _17585_/CLK _15875_/D vssd1 vssd1 vccd1 vccd1 _15875_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ _15004_/A _14826_/B vssd1 vssd1 vccd1 vccd1 _14826_/Y sky130_fd_sc_hd__nand2_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17614_ _17731_/CLK _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17545_ _18390_/CLK _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_1
X_14757_ hold3086/X _14772_/B _14756_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14757_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ hold2741/X _17147_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13708_ hold4209/X _13802_/B _13707_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17476_ _17478_/CLK _17476_/D vssd1 vssd1 vccd1 vccd1 _17476_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _15189_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16427_ _18370_/CLK _16427_/D vssd1 vssd1 vccd1 vccd1 _16427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13639_ hold5701/X _13829_/B _13638_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16358_ _18409_/CLK _16358_/D vssd1 vssd1 vccd1 vccd1 _16358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15309_ hold813/X _15485_/A2 _09392_/C hold610/X _15308_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5407 _16561_/Q vssd1 vssd1 vccd1 vccd1 hold5407/X sky130_fd_sc_hd__dlygate4sd3_1
X_16289_ _16311_/CLK _16289_/D vssd1 vssd1 vccd1 vccd1 _16289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5418 _11401_/X vssd1 vssd1 vccd1 vccd1 _16957_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5429 _16752_/Q vssd1 vssd1 vccd1 vccd1 hold5429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4706 _09661_/X vssd1 vssd1 vccd1 vccd1 _16377_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18028_ _18331_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4717 _16479_/Q vssd1 vssd1 vccd1 vccd1 hold4717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4728 _10216_/X vssd1 vssd1 vccd1 vccd1 _16562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4739 _16471_/Q vssd1 vssd1 vccd1 vccd1 hold4739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_395_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17867_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout206 _11207_/B vssd1 vssd1 vccd1 vccd1 _11789_/B sky130_fd_sc_hd__buf_4
Xfanout217 _10019_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__buf_4
X_09801_ _09918_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_324_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17207_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout228 _11095_/A2 vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__buf_4
XFILLER_0_227_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout239 _10477_/A2 vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__clkbuf_8
X_07993_ hold203/X _14681_/A vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09732_ _09933_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09663_ _09954_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ _09061_/A hold614/X vssd1 vssd1 vccd1 vccd1 _15929_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09594_ _10488_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08545_ _09061_/A hold280/X vssd1 vssd1 vccd1 vccd1 _15896_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _14529_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17814_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5930 _17549_/Q vssd1 vssd1 vccd1 vccd1 hold5930/X sky130_fd_sc_hd__dlygate4sd3_1
X_09028_ hold118/X hold429/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5941 _17553_/Q vssd1 vssd1 vccd1 vccd1 hold5941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5952 data_in[8] vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5963 data_in[21] vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5974 hold6031/X vssd1 vssd1 vccd1 vccd1 hold5974/X sky130_fd_sc_hd__buf_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5985 _15866_/Q vssd1 vssd1 vccd1 vccd1 hold5985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold29/X vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__clkbuf_4
Xhold5996 _18348_/Q vssd1 vssd1 vccd1 vccd1 hold5996/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__clkbuf_4
Xfanout751 fanout770/X vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout762 _13903_/A vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__buf_2
Xfanout773 fanout796/X vssd1 vssd1 vccd1 vccd1 _13750_/C1 sky130_fd_sc_hd__buf_4
X_13990_ _14330_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_176_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout784 _13941_/A vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__buf_4
Xfanout795 fanout796/X vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__clkbuf_4
X_12941_ hold3282/X _12940_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12942_/B sky130_fd_sc_hd__mux2_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15660_ _17236_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ hold3224/X _12871_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__mux2_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ hold1950/X _14610_/B _14610_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14611_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _13716_/A _11823_/B vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__or2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _17207_/CLK _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17330_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 _17330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14542_ hold2810/X _14541_/B _14541_/Y _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14542_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ hold4984/X _11658_/A _11753_/X vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ hold5130/X _11216_/B _10704_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17261_ _17261_/CLK _17261_/D vssd1 vssd1 vccd1 vccd1 _17261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _15099_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14473_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ _12219_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16212_ _17444_/CLK _16212_/D vssd1 vssd1 vccd1 vccd1 _16212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ hold2098/X hold3417/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13425_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ _11194_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _16702_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17192_ _18447_/CLK _17192_/D vssd1 vssd1 vccd1 vccd1 _17192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16143_ _16148_/CLK _16143_/D vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ hold1630/X hold3988/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10567_ _10603_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _16679_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12306_ hold4658/X _12213_/A _12305_/X vssd1 vssd1 vccd1 vccd1 _12306_/Y sky130_fd_sc_hd__a21oi_1
X_16074_ _17320_/CLK _16074_/D vssd1 vssd1 vccd1 vccd1 hold710/A sky130_fd_sc_hd__dfxtp_1
X_13286_ _13286_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ hold3714/X _10628_/B _10497_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10498_/X
+ sky130_fd_sc_hd__o211a_1
X_15025_ hold746/A _18296_/Q _15069_/S vssd1 vssd1 vccd1 vccd1 hold683/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12237_ _13773_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12168_ _13773_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or2_1
X_11119_ hold5056/X _11216_/B _11118_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12099_ _13797_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
X_16976_ _17851_/CLK _16976_/D vssd1 vssd1 vccd1 vccd1 _16976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput6 input6/A vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _17346_/CLK _15927_/D vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__dfxtp_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _17729_/CLK _15858_/D vssd1 vssd1 vccd1 vccd1 _15858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ hold2770/X _14828_/B _14808_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15789_ _17694_/CLK _15789_/D vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ hold2382/X _08336_/A2 _08329_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ _17534_/CLK _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ hold2674/X _08263_/A2 _08260_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17459_/CLK _17459_/D vssd1 vssd1 vccd1 vccd1 _17459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08192_ hold1992/X _08213_/B _08191_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5204 _16800_/Q vssd1 vssd1 vccd1 vccd1 hold5204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5215 _13603_/X vssd1 vssd1 vccd1 vccd1 _17654_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5226 _16480_/Q vssd1 vssd1 vccd1 vccd1 hold5226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5237 _10330_/X vssd1 vssd1 vccd1 vccd1 _16600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4503 hold5831/X vssd1 vssd1 vccd1 vccd1 hold5832/A sky130_fd_sc_hd__buf_4
Xhold5248 _17161_/Q vssd1 vssd1 vccd1 vccd1 hold5248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4514 _10918_/X vssd1 vssd1 vccd1 vccd1 _16796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5259 _12223_/X vssd1 vssd1 vccd1 vccd1 _17231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4525 _17710_/Q vssd1 vssd1 vccd1 vccd1 hold4525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4536 _09736_/X vssd1 vssd1 vccd1 vccd1 _16402_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3802 _16461_/Q vssd1 vssd1 vccd1 vccd1 hold3802/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4547 _17604_/Q vssd1 vssd1 vccd1 vccd1 hold4547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4558 _11128_/X vssd1 vssd1 vccd1 vccd1 _16866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3813 _11815_/X vssd1 vssd1 vccd1 vccd1 _17095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3824 _10522_/X vssd1 vssd1 vccd1 vccd1 _16664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4569 _17644_/Q vssd1 vssd1 vccd1 vccd1 hold4569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3835 _16362_/Q vssd1 vssd1 vccd1 vccd1 hold3835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3846 _12289_/X vssd1 vssd1 vccd1 vccd1 _17253_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3857 _15263_/X vssd1 vssd1 vccd1 vccd1 _15264_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3868 _16491_/Q vssd1 vssd1 vccd1 vccd1 hold3868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3879 _09895_/X vssd1 vssd1 vccd1 vccd1 _16455_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07976_ _15545_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ hold4181/X _10007_/B _09714_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09646_ hold4743/X _10049_/B _09645_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09646_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09577_ hold4855/X _10055_/B _09576_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09577_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08528_ hold215/X hold630/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold631/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08459_ hold2029/X _08488_/B _08458_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ hold5513/X _11762_/B _11469_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11470_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ hold2216/X hold3950/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_246_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18212_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13140_ hold4699/X _13139_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__mux2_1
X_10352_ hold1945/X _16608_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5760 _13723_/X vssd1 vssd1 vccd1 vccd1 _17694_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13071_ _13199_/A1 _13069_/X _13070_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13071_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5771 hold5926/X vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10283_ hold3116/X _16585_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__mux2_1
Xhold5782 hold5782/A vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_12
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5793 hold5936/X vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__dlygate4sd3_1
X_12022_ hold5218/X _12293_/B _12021_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16830_ _18063_/CLK _16830_/D vssd1 vssd1 vccd1 vccd1 _16830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout570 _07884_/Y vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__buf_6
Xfanout581 _13055_/X vssd1 vssd1 vccd1 vccd1 _13244_/S sky130_fd_sc_hd__buf_8
Xfanout592 _12970_/S vssd1 vssd1 vccd1 vccd1 _12748_/S sky130_fd_sc_hd__buf_4
X_16761_ _17994_/CLK _16761_/D vssd1 vssd1 vccd1 vccd1 _16761_/Q sky130_fd_sc_hd__dfxtp_1
X_13973_ hold1712/X _13995_/A2 _13972_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _13973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15712_ _17215_/CLK _15712_/D vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfxtp_1
X_12924_ _12996_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _17484_/D sky130_fd_sc_hd__and2_1
X_16692_ _18152_/CLK _16692_/D vssd1 vssd1 vccd1 vccd1 _16692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18431_ _18432_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15643_ _17153_/CLK _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _12921_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _17461_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11806_ hold4193/X _12031_/A2 _11805_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _11806_/X
+ sky130_fd_sc_hd__o211a_1
X_18362_ _18362_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ _17274_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12789_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _17438_/D sky130_fd_sc_hd__and2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17313_/CLK _17313_/D vssd1 vssd1 vccd1 vccd1 hold598/A sky130_fd_sc_hd__dfxtp_1
X_14525_ _14758_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _12310_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _17069_/D sky130_fd_sc_hd__nor2_1
X_18293_ _18293_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14456_ hold3234/X _14482_/A2 _14455_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14456_/X
+ sky130_fd_sc_hd__o211a_1
X_17244_ _17244_/CLK _17244_/D vssd1 vssd1 vccd1 vccd1 _17244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11668_ hold5441/X _11762_/B _11667_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11668_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13407_ _13779_/A _13407_/B vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__or2_1
X_10619_ _16697_/Q _10619_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17175_ _17207_/CLK _17175_/D vssd1 vssd1 vccd1 vccd1 _17175_/Q sky130_fd_sc_hd__dfxtp_1
X_14387_ _14782_/A hold2299/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11599_ hold5595/X _11768_/B _11598_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16126_ _16126_/CLK _16126_/D vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13338_ _13698_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16057_ _18407_/CLK _16057_/D vssd1 vssd1 vccd1 vccd1 _16057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ _13268_/X hold4619/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3109 _09085_/X vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15008_ hold972/X _15016_/B vssd1 vssd1 vccd1 vccd1 hold980/A sky130_fd_sc_hd__or2_1
Xhold2408 _14661_/X vssd1 vssd1 vccd1 vccd1 _18121_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2419 _09328_/X vssd1 vssd1 vccd1 vccd1 _16274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07830_ _14843_/A hold202/X vssd1 vssd1 vccd1 vccd1 _07871_/B sky130_fd_sc_hd__or2_4
Xhold1707 _08241_/X vssd1 vssd1 vccd1 vccd1 _15755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1718 _18207_/Q vssd1 vssd1 vccd1 vccd1 hold1718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 _17867_/Q vssd1 vssd1 vccd1 vccd1 hold1729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16959_ _17808_/CLK _16959_/D vssd1 vssd1 vccd1 vccd1 _16959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09500_ hold1875/X _16324_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _07785_/Y hold6004/X _15344_/A hold820/X vssd1 vssd1 vccd1 vccd1 hold821/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09362_ _09362_/A _09392_/B _09362_/C _09362_/D vssd1 vssd1 vccd1 vccd1 _09369_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08313_ _15537_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_176_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09293_ _15515_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08244_ _14517_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_33 fanout246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _14794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 hold525/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 hold915/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_77 _09339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_88 hold719/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08175_ _14164_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5001 _10345_/X vssd1 vssd1 vccd1 vccd1 _16605_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5012 _17063_/Q vssd1 vssd1 vccd1 vccd1 hold5012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5023 _12211_/X vssd1 vssd1 vccd1 vccd1 _17227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5034 _17083_/Q vssd1 vssd1 vccd1 vccd1 hold5034/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4300 _10957_/X vssd1 vssd1 vccd1 vccd1 _16809_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5045 _10939_/X vssd1 vssd1 vccd1 vccd1 _16803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5056 _16895_/Q vssd1 vssd1 vccd1 vccd1 hold5056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4311 _17036_/Q vssd1 vssd1 vccd1 vccd1 hold4311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5067 _10969_/X vssd1 vssd1 vccd1 vccd1 _16813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4322 _13456_/X vssd1 vssd1 vccd1 vccd1 _17605_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput140 hold990/X vssd1 vssd1 vccd1 vccd1 load_status[0] sky130_fd_sc_hd__buf_12
Xhold5078 _16759_/Q vssd1 vssd1 vccd1 vccd1 hold5078/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4333 _11413_/X vssd1 vssd1 vccd1 vccd1 _16961_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4344 _17680_/Q vssd1 vssd1 vccd1 vccd1 hold4344/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5089 _11524_/X vssd1 vssd1 vccd1 vccd1 _16998_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3610 _17380_/Q vssd1 vssd1 vccd1 vccd1 hold3610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4355 _11311_/X vssd1 vssd1 vccd1 vccd1 _16927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3621 _16511_/Q vssd1 vssd1 vccd1 vccd1 hold3621/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4366 _17737_/Q vssd1 vssd1 vccd1 vccd1 hold4366/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3632 _09565_/X vssd1 vssd1 vccd1 vccd1 _16345_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4377 _13666_/X vssd1 vssd1 vccd1 vccd1 _17675_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3643 _16676_/Q vssd1 vssd1 vccd1 vccd1 hold3643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4388 _10858_/X vssd1 vssd1 vccd1 vccd1 _16776_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3654 _09571_/X vssd1 vssd1 vccd1 vccd1 _16347_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4399 _16960_/Q vssd1 vssd1 vccd1 vccd1 hold4399/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3665 _11098_/X vssd1 vssd1 vccd1 vccd1 _16856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2920 _14480_/X vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2931 _18231_/Q vssd1 vssd1 vccd1 vccd1 hold2931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3676 _17418_/Q vssd1 vssd1 vccd1 vccd1 hold3676/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2942 _14635_/X vssd1 vssd1 vccd1 vccd1 _18108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3687 _16612_/Q vssd1 vssd1 vccd1 vccd1 hold3687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2953 _18120_/Q vssd1 vssd1 vccd1 vccd1 hold2953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3698 _13851_/Y vssd1 vssd1 vccd1 vccd1 _13852_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 _15100_/X vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2975 _14259_/X vssd1 vssd1 vccd1 vccd1 _17928_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07959_ hold2225/X _07991_/A2 _07958_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07959_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2986 _14081_/X vssd1 vssd1 vccd1 vccd1 _17843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2997 _18371_/Q vssd1 vssd1 vccd1 vccd1 hold2997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ hold1201/X _16814_/Q _11159_/C vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ hold2983/X _16367_/Q _10019_/C vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ hold1125/X hold3527/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12571_ hold2993/X _17368_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _15205_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_427_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17261_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11522_ hold1377/X hold3772/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__mux2_1
X_15290_ hold648/X _15486_/A2 _09357_/B hold339/X vssd1 vssd1 vccd1 vccd1 _15290_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ hold3185/X _14266_/B _14240_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _14241_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ hold2426/X hold4048/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10524_/A _10404_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__or2_1
X_14172_ _14403_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11384_ hold2494/X hold5569/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _13122_/X hold5912/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__mux2_1
X_10335_ _10554_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13054_/X
+ sky130_fd_sc_hd__and4b_4
Xhold5590 _10684_/X vssd1 vssd1 vccd1 vccd1 _16718_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17931_ _18055_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _10554_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ hold2987/X hold3774/X _12302_/C vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17862_ _17862_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
X_10197_ _10563_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16813_ _18014_/CLK _16813_/D vssd1 vssd1 vccd1 vccd1 _16813_/Q sky130_fd_sc_hd__dfxtp_1
X_17793_ _17825_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744_ _18006_/CLK _16744_/D vssd1 vssd1 vccd1 vccd1 _16744_/Q sky130_fd_sc_hd__dfxtp_1
X_13956_ _15517_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ hold2254/X hold3390/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_220_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16675_ _18231_/CLK _16675_/D vssd1 vssd1 vccd1 vccd1 _16675_/Q sky130_fd_sc_hd__dfxtp_1
X_13887_ hold3699/X _13779_/A _13886_/X vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18414_ _18422_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15626_ _17623_/CLK _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ hold2789/X hold3397/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__mux2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ _18377_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15557_ _15557_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__or2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ hold1181/X _17434_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14508_ hold1879/X _14535_/B _14507_/X _13903_/A vssd1 vssd1 vccd1 vccd1 _14508_/X
+ sky130_fd_sc_hd__o211a_1
X_15488_ hold563/X _15488_/A2 _15485_/X vssd1 vssd1 vccd1 vccd1 _15489_/D sky130_fd_sc_hd__a21o_1
X_18276_ _18276_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 input20/A vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_6
XFILLER_0_182_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _18428_/CLK _17227_/D vssd1 vssd1 vccd1 vccd1 _17227_/Q sky130_fd_sc_hd__dfxtp_1
Xinput31 hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14439_ _15173_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 input42/A vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput53 input53/A vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_4
XFILLER_0_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput64 input64/A vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_6
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _17189_/CLK _17158_/D vssd1 vssd1 vccd1 vccd1 _17158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold815 hold815/A vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 hold837/A vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16109_ _17332_/CLK _16109_/D vssd1 vssd1 vccd1 vccd1 hold592/A sky130_fd_sc_hd__dfxtp_1
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ hold2695/X hold5280/X _11159_/C vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17089_ _17871_/CLK _17089_/D vssd1 vssd1 vccd1 vccd1 _17089_/Q sky130_fd_sc_hd__dfxtp_1
Xhold859 hold859/A vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ _15344_/A hold898/X vssd1 vssd1 vccd1 vccd1 _16083_/D sky130_fd_sc_hd__and2_1
XFILLER_0_228_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2205 _16239_/Q vssd1 vssd1 vccd1 vccd1 hold2205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2216 _18187_/Q vssd1 vssd1 vccd1 vccd1 hold2216/X sky130_fd_sc_hd__dlygate4sd3_1
X_08862_ hold292/X hold799/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold800/A sky130_fd_sc_hd__mux2_1
Xhold2227 _15671_/Q vssd1 vssd1 vccd1 vccd1 hold2227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2238 _18350_/Q vssd1 vssd1 vccd1 vccd1 hold2238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 _14283_/X vssd1 vssd1 vccd1 vccd1 _17940_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _07844_/X vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 _15771_/Q vssd1 vssd1 vccd1 vccd1 hold1515/X sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ _15531_/A _14988_/A hold944/X _14984_/A vssd1 vssd1 vccd1 vccd1 _07813_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1526 _13944_/X vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08793_ hold150/X hold176/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__mux2_1
Xhold1537 _08390_/X vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 _09302_/X vssd1 vssd1 vccd1 vccd1 _16261_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1559 _15800_/Q vssd1 vssd1 vccd1 vccd1 hold1559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09414_ _09438_/B _16293_/Q vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09345_ _15555_/A _15173_/A _15551_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09359_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_176_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _12759_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _16249_/D sky130_fd_sc_hd__and2_1
XFILLER_0_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08227_ hold689/A hold764/A hold732/A hold752/A vssd1 vssd1 vccd1 vccd1 _15128_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_106_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ _15509_/A hold1163/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ hold2612/X _08088_/B _08088_/Y _08127_/A vssd1 vssd1 vccd1 vccd1 _08089_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4130 _13522_/X vssd1 vssd1 vccd1 vccd1 _17627_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10120_ hold5260/X _10598_/B _10119_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _10120_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4141 _17615_/Q vssd1 vssd1 vccd1 vccd1 hold4141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4152 _12184_/X vssd1 vssd1 vccd1 vccd1 _17218_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4163 _10285_/X vssd1 vssd1 vccd1 vccd1 _16585_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4174 _11884_/X vssd1 vssd1 vccd1 vccd1 _17118_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3440 _17269_/Q vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4185 _17706_/Q vssd1 vssd1 vccd1 vccd1 hold4185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10051_ _10603_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _16507_/D sky130_fd_sc_hd__nor2_1
Xhold4196 _10468_/X vssd1 vssd1 vccd1 vccd1 _16646_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3451 _12073_/X vssd1 vssd1 vccd1 vccd1 _17181_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3462 _17653_/Q vssd1 vssd1 vccd1 vccd1 hold3462/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3473 _12566_/X vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3484 _17611_/Q vssd1 vssd1 vccd1 vccd1 hold3484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2750 _18111_/Q vssd1 vssd1 vccd1 vccd1 hold2750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3495 _11986_/X vssd1 vssd1 vccd1 vccd1 _17152_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2761 _15746_/Q vssd1 vssd1 vccd1 vccd1 hold2761/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2772 _15747_/Q vssd1 vssd1 vccd1 vccd1 hold2772/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2783 _15534_/X vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2794 _07903_/X vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13825_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _17723_/D sky130_fd_sc_hd__nor2_1
X_14790_ _15183_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__or2_1
XFILLER_0_199_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ hold4541/X _13856_/B _13740_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _11052_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16460_ _18371_/CLK _16460_/D vssd1 vssd1 vccd1 vccd1 _16460_/Q sky130_fd_sc_hd__dfxtp_1
X_13672_ hold5691/X _13817_/B _13671_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _13672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ _11643_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _16305_/Q _15477_/A2 _15487_/B1 hold283/X _15410_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/D sky130_fd_sc_hd__a221o_1
X_12623_ hold3310/X _12622_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12623_/X sky130_fd_sc_hd__mux2_1
X_16391_ _18276_/CLK _16391_/D vssd1 vssd1 vccd1 vccd1 _16391_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _15489_/A _15342_/B _15342_/C _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/X
+ sky130_fd_sc_hd__or4_1
X_18130_ _18208_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_261_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18067_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12554_ hold3595/X _12553_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _11706_/A _11505_/B vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__or2_1
X_15273_ _15490_/A1 _15265_/X _15272_/X _15490_/B1 hold5842/A vssd1 vssd1 vccd1 vccd1
+ _15273_/X sky130_fd_sc_hd__a32o_1
X_18061_ _18061_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
X_12485_ hold44/X _12445_/A _12445_/B _12484_/X _12444_/A vssd1 vssd1 vccd1 vccd1
+ hold45/A sky130_fd_sc_hd__o311a_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14224_ _14974_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__or2_1
X_17012_ _17858_/CLK _17012_/D vssd1 vssd1 vccd1 vccd1 _17012_/Q sky130_fd_sc_hd__dfxtp_1
X_11436_ _11631_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14155_ hold2707/X _14148_/B _14154_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _14155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ _11643_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _17564_/Q _17098_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10318_ hold4889/X _10649_/B _10317_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14086_ _15539_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__or2_1
X_11298_ _12285_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__or2_1
X_13037_ _13037_/A hold961/X vssd1 vssd1 vccd1 vccd1 _17522_/D sky130_fd_sc_hd__and2_1
X_17914_ _18006_/CLK _17914_/D vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_1
X_10249_ hold4970/X _10631_/B _10248_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ _17877_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _17808_/CLK _17776_/D vssd1 vssd1 vccd1 vccd1 _17776_/Q sky130_fd_sc_hd__dfxtp_1
X_14988_ _14988_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16727_ _18124_/CLK _16727_/D vssd1 vssd1 vccd1 vccd1 _16727_/Q sky130_fd_sc_hd__dfxtp_1
X_13939_ _13943_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _17775_/D sky130_fd_sc_hd__and2_1
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_349_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17681_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16658_ _18214_/CLK _16658_/D vssd1 vssd1 vccd1 vccd1 _16658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15609_ _17257_/CLK _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16589_ _18209_/CLK _16589_/D vssd1 vssd1 vccd1 vccd1 _16589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09130_ _15513_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__or2_1
X_18328_ _18360_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09061_ _09061_/A hold542/X vssd1 vssd1 vccd1 vccd1 _16147_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18259_ _18387_/CLK hold987/X vssd1 vssd1 vccd1 vccd1 hold986/A sky130_fd_sc_hd__dfxtp_1
X_08012_ hold2987/X _08029_/B _08011_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _08012_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 hold807/X vssd1 vssd1 vccd1 vccd1 hold808/A sky130_fd_sc_hd__buf_6
Xhold612 hold612/A vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold623 hold623/A vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold634 hold634/A vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold645 hold645/A vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 hold656/A vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold667 hold667/A vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold678 hold678/A vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__or2_1
Xhold689 hold689/A vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_65_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18044_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2002 _18201_/Q vssd1 vssd1 vccd1 vccd1 hold2002/X sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ hold607/X hold836/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold837/A sky130_fd_sc_hd__mux2_1
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2013 _07812_/Y vssd1 vssd1 vccd1 vccd1 hold2013/X sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ _09933_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__or2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _14145_/X vssd1 vssd1 vccd1 vccd1 _17874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2035 _16193_/Q vssd1 vssd1 vccd1 vccd1 hold2035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2046 _07808_/X vssd1 vssd1 vccd1 vccd1 _17752_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 hold1402/X vssd1 vssd1 vccd1 vccd1 hold1301/X sky130_fd_sc_hd__buf_1
XFILLER_0_97_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08845_ _12408_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _16041_/D sky130_fd_sc_hd__and2_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 _08514_/X vssd1 vssd1 vccd1 vccd1 _15884_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 hold6037/X vssd1 vssd1 vccd1 vccd1 hold1312/X sky130_fd_sc_hd__buf_1
Xhold1323 hold6023/X vssd1 vssd1 vccd1 vccd1 _09447_/C sky130_fd_sc_hd__clkbuf_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2068 _17848_/Q vssd1 vssd1 vccd1 vccd1 hold2068/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 _15848_/Q vssd1 vssd1 vccd1 vccd1 hold2079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 hold1440/X vssd1 vssd1 vccd1 vccd1 hold1334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 _14793_/X vssd1 vssd1 vccd1 vccd1 _18184_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1356 hold1356/A vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__buf_12
XFILLER_0_225_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08776_ _15394_/A hold608/X vssd1 vssd1 vccd1 vccd1 _16008_/D sky130_fd_sc_hd__and2_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1367 _15574_/Q vssd1 vssd1 vccd1 vccd1 hold1367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 _14083_/X vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1389 _18236_/Q vssd1 vssd1 vccd1 vccd1 hold1389/X sky130_fd_sc_hd__buf_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09328_ hold2418/X _09325_/B _09327_/X _12600_/A vssd1 vssd1 vccd1 vccd1 _09328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _15535_/A hold1196/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ _12273_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _12340_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _16897_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11152_ _12310_/A _11152_/B vssd1 vssd1 vccd1 vccd1 _16874_/D sky130_fd_sc_hd__nor2_1
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ hold1899/X hold4627/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ _17322_/CLK _15960_/D vssd1 vssd1 vccd1 vccd1 hold456/A sky130_fd_sc_hd__dfxtp_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ hold4715/X _11177_/B _11082_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _11083_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3270 _17492_/Q vssd1 vssd1 vccd1 vccd1 hold3270/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10034_ _16502_/Q _10034_/B _10034_/C vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__and3_1
X_14911_ hold2480/X _14896_/Y _14910_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14911_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3281 _17354_/Q vssd1 vssd1 vccd1 vccd1 hold3281/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3292 _17381_/Q vssd1 vssd1 vccd1 vccd1 hold3292/X sky130_fd_sc_hd__dlygate4sd3_1
X_15891_ _17339_/CLK _15891_/D vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__dfxtp_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2580 _09217_/X vssd1 vssd1 vccd1 vccd1 _16220_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _17726_/CLK _17630_/D vssd1 vssd1 vccd1 vccd1 _17630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _14843_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14842_/Y sky130_fd_sc_hd__nor2_2
Xhold2591 _07933_/X vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 hold1890/A vssd1 vssd1 vccd1 vccd1 input67/A sky130_fd_sc_hd__dlygate4sd3_1
X_17561_ _17721_/CLK _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
X_14773_ hold1990/X _14772_/B _14772_/Y _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14773_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _13782_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16512_ _18108_/CLK _16512_/D vssd1 vssd1 vccd1 vccd1 _16512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_442_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17722_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13724_ hold1164/X hold5713/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10936_ hold4553/X _11789_/B _10935_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _10936_/X
+ sky130_fd_sc_hd__o211a_1
X_17492_ _17509_/CLK _17492_/D vssd1 vssd1 vccd1 vccd1 _17492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16443_ _18322_/CLK _16443_/D vssd1 vssd1 vccd1 vccd1 _16443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ hold5471/X _10019_/B _10866_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10867_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13655_ hold2445/X hold3531/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ _12606_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _17378_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _18349_/CLK _16374_/D vssd1 vssd1 vccd1 vccd1 _16374_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ hold2300/X hold3482/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__mux2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ hold4753/X _11177_/B _10797_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18113_ _18113_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15325_ _15325_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15325_/X sky130_fd_sc_hd__or2_1
X_12537_ _12606_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _17355_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18044_ _18044_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15256_ _17329_/Q _15448_/B1 _15485_/B1 hold462/X vssd1 vssd1 vccd1 vccd1 _15256_/X
+ sky130_fd_sc_hd__a22o_1
X_12468_ _17327_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14207_ hold1654/X _14202_/B _14206_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14207_/X
+ sky130_fd_sc_hd__o211a_1
X_11419_ hold4439/X _11801_/B _11418_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11419_/X
+ sky130_fd_sc_hd__o211a_1
X_15187_ hold746/X _15211_/B vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__or2_1
X_12399_ hold163/X hold320/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14138_ _15211_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ hold2293/X _14107_/A2 _14068_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _12386_/A hold589/X vssd1 vssd1 vccd1 vccd1 _15937_/D sky130_fd_sc_hd__and2_1
X_17828_ _17860_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08561_ _09053_/A hold119/X vssd1 vssd1 vccd1 vccd1 _15904_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _17887_/CLK _17759_/D vssd1 vssd1 vccd1 vccd1 _17759_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_183_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18391_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08492_ _14330_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17340_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ hold2502/X _09119_/A2 _09112_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ hold607/X hold637/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold638/A sky130_fd_sc_hd__mux2_1
Xhold420 hold420/A vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/A vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold453 input9/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold464 hold464/A vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 hold524/X vssd1 vssd1 vccd1 vccd1 hold525/A sky130_fd_sc_hd__buf_6
XFILLER_0_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout900 hold746/X vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__clkbuf_16
Xhold497 input28/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__buf_1
XFILLER_0_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout911 hold1079/X vssd1 vssd1 vccd1 vccd1 hold1080/A sky130_fd_sc_hd__buf_6
XFILLER_0_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout922 hold971/X vssd1 vssd1 vccd1 vccd1 hold972/A sky130_fd_sc_hd__buf_4
X_09946_ hold5673/X _10070_/B _09945_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09946_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout933 hold1015/X vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout944 hold1301/X vssd1 vssd1 vccd1 vccd1 hold1302/A sky130_fd_sc_hd__buf_6
XFILLER_0_216_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ hold3681/X _10565_/B _09876_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09877_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _13951_/X vssd1 vssd1 vccd1 vccd1 _17780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _08190_/X vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 input51/X vssd1 vssd1 vccd1 vccd1 hold1142/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ hold271/X hold370/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__mux2_1
Xhold1153 _15493_/X vssd1 vssd1 vccd1 vccd1 _15494_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _15724_/Q vssd1 vssd1 vccd1 vccd1 hold1164/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1175 _14877_/X vssd1 vssd1 vccd1 vccd1 _18225_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1186 _15689_/Q vssd1 vssd1 vccd1 vccd1 hold1186/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ hold118/X hold814/X _08759_/S vssd1 vssd1 vccd1 vccd1 hold815/A sky130_fd_sc_hd__mux2_1
Xhold1197 _17516_/Q vssd1 vssd1 vccd1 vccd1 hold1197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _12367_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _17080_/D sky130_fd_sc_hd__nor2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10721_ hold2351/X hold4960/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _13767_/A _13440_/B vssd1 vssd1 vccd1 vccd1 _13440_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10652_ hold1939/X hold4155/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _13791_/A _13371_/B vssd1 vssd1 vccd1 vccd1 _13371_/X sky130_fd_sc_hd__or2_1
X_10583_ _16685_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__and3_1
XFILLER_0_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15110_ hold988/X _15113_/B _15109_/Y _15044_/A vssd1 vssd1 vccd1 vccd1 hold989/A
+ sky130_fd_sc_hd__o211a_1
X_12322_ _13825_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _17264_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16090_ _17306_/CLK _16090_/D vssd1 vssd1 vccd1 vccd1 hold739/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ _14988_/A hold2799/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__mux2_1
X_12253_ _12347_/A _12347_/B _12252_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11204_ _16892_/Q _11753_/B _11204_/C vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__and3_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ hold4151/X _12374_/B _12183_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _12184_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ hold1960/X _16869_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _11136_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ _17891_/CLK _16992_/D vssd1 vssd1 vccd1 vccd1 _16992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15943_ _18415_/CLK _15943_/D vssd1 vssd1 vccd1 vccd1 _15943_/Q sky130_fd_sc_hd__dfxtp_1
X_11066_ hold1416/X hold5180/X _11201_/C vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__mux2_1
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _13158_/A _09963_/A _10016_/X vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _17585_/CLK _15874_/D vssd1 vssd1 vccd1 vccd1 _15874_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _17613_/CLK _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ hold2115/X _14828_/B _14824_/Y _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14825_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _18390_/CLK _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _14988_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11968_ hold3456/X _12347_/B _11967_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _13713_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__or2_1
X_17475_ _17478_/CLK _17475_/D vssd1 vssd1 vccd1 vccd1 _17475_/Q sky130_fd_sc_hd__dfxtp_1
X_10919_ hold2094/X _16797_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14687_ hold1912/X _14720_/B _14686_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14687_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11899_ hold4342/X _13877_/B _11898_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ _18395_/CLK _16426_/D vssd1 vssd1 vccd1 vccd1 _16426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13638_ _13734_/A _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16357_ _18300_/CLK _16357_/D vssd1 vssd1 vccd1 vccd1 _16357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ _13746_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13569_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15308_ hold838/X _09386_/A _15451_/A2 hold778/X vssd1 vssd1 vccd1 vccd1 _15308_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5408 _10117_/X vssd1 vssd1 vccd1 vccd1 _16529_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16288_ _16312_/CLK _16288_/D vssd1 vssd1 vccd1 vccd1 _16288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5419 _17166_/Q vssd1 vssd1 vccd1 vccd1 hold5419/X sky130_fd_sc_hd__dlygate4sd3_1
X_18027_ _18032_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
X_15239_ hold649/X _15485_/A2 _15488_/A2 hold786/X _15238_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_125_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4707 _16736_/Q vssd1 vssd1 vccd1 vccd1 hold4707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4718 _09871_/X vssd1 vssd1 vccd1 vccd1 _16447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4729 _17115_/Q vssd1 vssd1 vccd1 vccd1 hold4729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09800_ hold2755/X _16424_/Q _10019_/C vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__mux2_1
Xfanout207 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__buf_4
Xfanout218 _10025_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout229 fanout246/X vssd1 vssd1 vccd1 vccd1 _11095_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07992_ hold764/A hold732/X hold752/X hold689/X vssd1 vssd1 vccd1 vccd1 _14681_/A
+ sky130_fd_sc_hd__nand4b_4
XFILLER_0_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09731_ _18312_/Q hold4000/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09662_ hold1342/X hold4735/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_364_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08613_ hold596/X hold613/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold614/A sky130_fd_sc_hd__mux2_1
X_09593_ hold1702/X _13310_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08544_ hold47/X _15896_/Q _08592_/S vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__mux2_1
XFILLER_0_167_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ hold5985/X _08486_/B _08474_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08475_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_6_9_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_80_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09027_ _15364_/A hold675/X vssd1 vssd1 vccd1 vccd1 _16130_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5920 _16925_/Q vssd1 vssd1 vccd1 vccd1 hold5920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5931 _17534_/Q vssd1 vssd1 vccd1 vccd1 hold5931/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5942 _17533_/Q vssd1 vssd1 vccd1 vccd1 hold5942/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5953 data_in[1] vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5964 data_in[19] vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 input30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold261 hold61/X vssd1 vssd1 vccd1 vccd1 input20/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5975 _15760_/Q vssd1 vssd1 vccd1 vccd1 hold5975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5986 data_in[27] vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5997 _18274_/Q vssd1 vssd1 vccd1 vccd1 hold5997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout730 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__buf_4
Xfanout741 _15454_/A vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__buf_4
X_09929_ hold1054/X _16467_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__mux2_1
Xfanout752 fanout770/X vssd1 vssd1 vccd1 vccd1 _13777_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_205_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout763 fanout770/X vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__buf_4
Xfanout774 _08125_/A vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__buf_4
Xfanout785 fanout796/X vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout796 fanout847/X vssd1 vssd1 vccd1 vccd1 fanout796/X sky130_fd_sc_hd__buf_4
XFILLER_0_198_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12940_ hold1063/X hold3280/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ hold3039/X hold3149/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12871_/X sky130_fd_sc_hd__mux2_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _15004_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__nand2_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11822_ hold2074/X hold3569/X _12302_/C vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _17145_/CLK _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14541_ _14774_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__nand2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _17075_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__and3_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11094_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__or2_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17260_ _17260_/CLK _17260_/D vssd1 vssd1 vccd1 vccd1 _17260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ hold2737/X _17052_/Q _12314_/C vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__mux2_1
X_14472_ hold2634/X _14482_/A2 _14471_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14472_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _18438_/CLK hold992/X vssd1 vssd1 vccd1 vccd1 hold991/A sky130_fd_sc_hd__dfxtp_1
X_10635_ hold4619/X _11100_/A _10634_/X vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13423_ hold4010/X _13802_/B _13422_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17191_ _17194_/CLK _17191_/D vssd1 vssd1 vccd1 vccd1 _17191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16142_ _17339_/CLK _16142_/D vssd1 vssd1 vccd1 vccd1 hold489/A sky130_fd_sc_hd__dfxtp_1
X_13354_ hold5735/X _13832_/B _13353_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _13354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ hold3543/X _10560_/A _10565_/X vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _17259_/Q _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12305_/X sky130_fd_sc_hd__and3_1
XFILLER_0_87_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16073_ _17320_/CLK _16073_/D vssd1 vssd1 vccd1 vccd1 hold758/A sky130_fd_sc_hd__dfxtp_1
X_13285_ _13284_/X hold3571/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15024_ _15024_/A _15024_/B vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__and2_1
X_12236_ hold1350/X _17236_/Q _13868_/C vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12167_ hold2605/X hold3450/X _12251_/S vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11118_ _11121_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12098_ hold1294/X _17190_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__mux2_1
X_16975_ _17821_/CLK _16975_/D vssd1 vssd1 vccd1 vccd1 _16975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ _16077_/CLK _15926_/D vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _11052_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _17731_/CLK _15857_/D vssd1 vssd1 vccd1 vccd1 _15857_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _14862_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__or2_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _17693_/CLK _15788_/D vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17527_ _17534_/CLK _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_1
X_14739_ hold1338/X _14774_/B _14738_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14739_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08260_ _15539_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _17459_/CLK _17458_/D vssd1 vssd1 vccd1 vccd1 _17458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _18384_/CLK _16409_/D vssd1 vssd1 vccd1 vccd1 _16409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08191_ _15199_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _18452_/CLK _17389_/D vssd1 vssd1 vccd1 vccd1 _17389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5205 _10834_/X vssd1 vssd1 vccd1 vccd1 _16768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5216 _17032_/Q vssd1 vssd1 vccd1 vccd1 hold5216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5227 _09874_/X vssd1 vssd1 vccd1 vccd1 _16448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5238 _17718_/Q vssd1 vssd1 vccd1 vccd1 hold5238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4504 _15303_/X vssd1 vssd1 vccd1 vccd1 _15304_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5249 _11917_/X vssd1 vssd1 vccd1 vccd1 _17129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4515 _17090_/Q vssd1 vssd1 vccd1 vccd1 hold4515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4526 _13675_/X vssd1 vssd1 vccd1 vccd1 _17678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4537 _16897_/Q vssd1 vssd1 vccd1 vccd1 hold4537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3803 _09817_/X vssd1 vssd1 vccd1 vccd1 _16429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4548 _13357_/X vssd1 vssd1 vccd1 vccd1 _17572_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3814 _17410_/Q vssd1 vssd1 vccd1 vccd1 hold3814/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4559 _17668_/Q vssd1 vssd1 vccd1 vccd1 hold4559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3825 _17112_/Q vssd1 vssd1 vccd1 vccd1 hold3825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3836 _09520_/X vssd1 vssd1 vccd1 vccd1 _16330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3847 _17401_/Q vssd1 vssd1 vccd1 vccd1 hold3847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3858 _16437_/Q vssd1 vssd1 vccd1 vccd1 hold3858/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3869 _09907_/X vssd1 vssd1 vccd1 vccd1 _16459_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07975_ hold2015/X _07978_/B _07974_/Y _08353_/A vssd1 vssd1 vccd1 vccd1 _07975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09714_ _09936_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09645_ _09954_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ _09960_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__or2_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _15491_/A hold726/X vssd1 vssd1 vccd1 vccd1 _15888_/D sky130_fd_sc_hd__and2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _15517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _15826_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ hold4053/X _10628_/B _10419_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10420_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10351_ hold4974/X _10631_/B _10350_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ _13070_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__or2_1
Xhold5750 _13768_/X vssd1 vssd1 vccd1 vccd1 _17709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10282_ hold4757/X _10571_/B _10281_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10282_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5761 _17632_/Q vssd1 vssd1 vccd1 vccd1 hold5761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5772 output90/X vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_12
Xhold5783 hold5931/X vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12021_ _12288_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__or2_1
Xhold5794 output80/X vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_286_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_215_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_206_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout560 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08097_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_205_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 _07871_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__buf_8
XFILLER_0_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout582 _13055_/X vssd1 vssd1 vccd1 vccd1 _13308_/S sky130_fd_sc_hd__buf_8
X_16760_ _18200_/CLK _16760_/D vssd1 vssd1 vccd1 vccd1 _16760_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout593 _12826_/S vssd1 vssd1 vccd1 vccd1 _12808_/S sky130_fd_sc_hd__buf_6
X_13972_ _15207_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15711_ _17903_/CLK _15711_/D vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfxtp_1
X_12923_ hold3294/X _12922_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12924_/B sky130_fd_sc_hd__mux2_1
X_16691_ _18215_/CLK _16691_/D vssd1 vssd1 vccd1 vccd1 _16691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ _18430_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15642_ _17237_/CLK _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ hold3304/X _12853_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_201_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18361_ _18387_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_11805_ _12024_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__or2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _17171_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12785_ hold3308/X _12784_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__mux2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17312_ _17332_/CLK _17312_/D vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14524_ hold3088/X _14541_/B _14523_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14524_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18292_/CLK hold721/X vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ hold4674/X _11643_/A _11735_/X vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17243_ _17590_/CLK _17243_/D vssd1 vssd1 vccd1 vccd1 _17243_/Q sky130_fd_sc_hd__dfxtp_1
X_14455_ _15189_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11667_ _11667_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13406_ hold1289/X _17589_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13407_/B sky130_fd_sc_hd__mux2_1
X_10618_ _11194_/A _10618_/B vssd1 vssd1 vccd1 vccd1 _16696_/D sky130_fd_sc_hd__nor2_1
X_17174_ _17270_/CLK _17174_/D vssd1 vssd1 vccd1 vccd1 _17174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14386_ _14386_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__and2_1
X_11598_ _11694_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _17326_/CLK _16125_/D vssd1 vssd1 vccd1 vccd1 hold543/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10549_ hold3952/X _10646_/B _10548_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10549_/X
+ sky130_fd_sc_hd__o211a_1
X_13337_ hold1061/X hold4643/X _13817_/C vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _18410_/CLK _16056_/D vssd1 vssd1 vccd1 vccd1 hold536/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ hold4929/X _13267_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ hold1043/X hold514/X _15006_/Y _15007_/C1 vssd1 vssd1 vccd1 vccd1 _15007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12219_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _13199_/A1 _13197_/X _13198_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2409 _17842_/Q vssd1 vssd1 vccd1 vccd1 hold2409/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1708 _17836_/Q vssd1 vssd1 vccd1 vccd1 hold1708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 _14839_/X vssd1 vssd1 vccd1 vccd1 _18207_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16958_ _17804_/CLK _16958_/D vssd1 vssd1 vccd1 vccd1 _16958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ _16089_/CLK _15909_/D vssd1 vssd1 vccd1 vccd1 hold634/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16889_ _17999_/CLK _16889_/D vssd1 vssd1 vccd1 vccd1 _16889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09430_ hold819/X _16301_/Q vssd1 vssd1 vccd1 vccd1 hold820/A sky130_fd_sc_hd__or2_1
XFILLER_0_232_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ _09366_/A _09364_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ hold1462/X _08323_/B _08311_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _08312_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ hold1583/X _09338_/A2 _09291_/X _12606_/A vssd1 vssd1 vccd1 vccd1 _09292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ hold2077/X _08263_/A2 _08242_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _14862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_56 hold607/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_67 hold954/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08174_ hold203/X _15182_/A vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__or2_4
XANTENNA_78 hold5856/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 hold719/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5002 _16900_/Q vssd1 vssd1 vccd1 vccd1 hold5002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5013 _11623_/X vssd1 vssd1 vccd1 vccd1 _17031_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5024 _17132_/Q vssd1 vssd1 vccd1 vccd1 hold5024/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5035 _11683_/X vssd1 vssd1 vccd1 vccd1 _17051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4301 _17215_/Q vssd1 vssd1 vccd1 vccd1 hold4301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5046 _16753_/Q vssd1 vssd1 vccd1 vccd1 hold5046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5057 _11119_/X vssd1 vssd1 vccd1 vccd1 _16863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4312 _11542_/X vssd1 vssd1 vccd1 vccd1 _17004_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4323 _17639_/Q vssd1 vssd1 vccd1 vccd1 hold4323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput130 hold5884/X vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_12
XFILLER_0_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5068 _16919_/Q vssd1 vssd1 vccd1 vccd1 hold5068/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput141 _13043_/C vssd1 vssd1 vccd1 vccd1 load_status[1] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5079 _10711_/X vssd1 vssd1 vccd1 vccd1 _16727_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4334 _17619_/Q vssd1 vssd1 vccd1 vccd1 hold4334/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4345 _13585_/X vssd1 vssd1 vccd1 vccd1 _17648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3600 _16907_/Q vssd1 vssd1 vccd1 vccd1 hold3600/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4356 _17609_/Q vssd1 vssd1 vccd1 vccd1 hold4356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3611 _17108_/Q vssd1 vssd1 vccd1 vccd1 hold3611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3622 _09967_/X vssd1 vssd1 vccd1 vccd1 _16479_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4367 _13756_/X vssd1 vssd1 vccd1 vccd1 _17705_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3633 hold4107/X vssd1 vssd1 vccd1 vccd1 _13814_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4378 _17057_/Q vssd1 vssd1 vccd1 vccd1 hold4378/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3644 _10462_/X vssd1 vssd1 vccd1 vccd1 _16644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4389 _17617_/Q vssd1 vssd1 vccd1 vccd1 hold4389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3655 _16475_/Q vssd1 vssd1 vccd1 vccd1 hold3655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2910 _14534_/X vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3666 hold4384/X vssd1 vssd1 vccd1 vccd1 _13838_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2921 _17952_/Q vssd1 vssd1 vccd1 vccd1 hold2921/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3677 _16571_/Q vssd1 vssd1 vccd1 vccd1 hold3677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2932 _14889_/X vssd1 vssd1 vccd1 vccd1 _18231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3688 _10270_/X vssd1 vssd1 vccd1 vccd1 _16580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 _18069_/Q vssd1 vssd1 vccd1 vccd1 hold2943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2954 _14659_/X vssd1 vssd1 vccd1 vccd1 _18120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3699 _17589_/Q vssd1 vssd1 vccd1 vccd1 hold3699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2965 _15699_/Q vssd1 vssd1 vccd1 vccd1 hold2965/X sky130_fd_sc_hd__dlygate4sd3_1
X_07958_ _14862_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07958_/X sky130_fd_sc_hd__or2_1
Xhold2976 _15675_/Q vssd1 vssd1 vccd1 vccd1 hold2976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2987 _15647_/Q vssd1 vssd1 vccd1 vccd1 hold2987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 _15180_/X vssd1 vssd1 vccd1 vccd1 _18371_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07889_ hold1256/X _07924_/B _07888_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _07889_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ hold5350/X _10034_/B _09627_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09559_ hold3619/X _10037_/B _09558_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09559_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ _12960_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _17366_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ hold3746/X _11617_/A2 _11520_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11521_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _15189_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__or2_1
X_11452_ hold5222/X _11738_/B _11451_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ hold1555/X hold4938/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10404_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14171_ hold2911/X _14198_/B _14170_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11383_ hold5637/X _11789_/B _11382_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10334_ hold1338/X _16602_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _17566_/Q _17100_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_239_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13053_ _13053_/A _13056_/C _13055_/C _17523_/Q vssd1 vssd1 vccd1 vccd1 _13053_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_221_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5580 _11062_/X vssd1 vssd1 vccd1 vccd1 _16844_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17930_ _18063_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10265_ hold2380/X _16579_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__mux2_1
Xhold5591 _16776_/Q vssd1 vssd1 vccd1 vccd1 hold5591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12004_ hold5346/X _13798_/A2 _12003_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12004_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4890 _10318_/X vssd1 vssd1 vccd1 vccd1 _16596_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17861_ _17902_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
X_10196_ hold1771/X _16556_/Q _10580_/C vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16812_ _18459_/CLK _16812_/D vssd1 vssd1 vccd1 vccd1 _16812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _17884_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout390 _14626_/Y vssd1 vssd1 vccd1 vccd1 _14666_/B sky130_fd_sc_hd__buf_6
XFILLER_0_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16743_ _18010_/CLK _16743_/D vssd1 vssd1 vccd1 vccd1 _16743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13955_ hold2856/X _13995_/A2 _13954_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _13955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12909_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _17478_/D sky130_fd_sc_hd__and2_1
X_16674_ _18166_/CLK _16674_/D vssd1 vssd1 vccd1 vccd1 _16674_/Q sky130_fd_sc_hd__dfxtp_1
X_13886_ _17749_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__and3_1
X_18413_ _18413_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
X_15625_ _17189_/CLK _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12837_ _12870_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _17455_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18386_/CLK hold736/X vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15556_ hold2913/X _15560_/A2 _15555_/X _12759_/A vssd1 vssd1 vccd1 vccd1 _15556_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12768_ _12768_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _17432_/D sky130_fd_sc_hd__and2_1
XFILLER_0_33_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ _14794_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14507_/X sky130_fd_sc_hd__or2_1
X_18275_ _18349_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _12310_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _17063_/D sky130_fd_sc_hd__nor2_1
X_15487_ _17324_/Q _15487_/A2 _15487_/B1 hold302/X _15486_/X vssd1 vssd1 vccd1 vccd1
+ _15489_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12699_ _12768_/A _12699_/B vssd1 vssd1 vccd1 vccd1 _17409_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17226_ _17258_/CLK _17226_/D vssd1 vssd1 vccd1 vccd1 _17226_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 input10/A vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
X_14438_ hold1201/X _14446_/A2 _14437_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 input21/A vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_6
Xinput32 input32/A vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput43 input43/A vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 input54/A vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_6
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17157_ _17157_/CLK _17157_/D vssd1 vssd1 vccd1 vccd1 _17157_/Q sky130_fd_sc_hd__dfxtp_1
X_14369_ _15103_/A hold2823/X hold333/X vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
Xhold805 la_data_in[25] vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_137_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16127_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16108_ _17335_/CLK _16108_/D vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
Xhold827 hold827/A vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 hold838/A vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 hold849/A vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _17870_/CLK _17088_/D vssd1 vssd1 vccd1 vccd1 _17088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16039_ _17298_/CLK _16039_/D vssd1 vssd1 vccd1 vccd1 hold878/A sky130_fd_sc_hd__dfxtp_1
X_08930_ hold498/X hold897/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold898/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2206 _16258_/Q vssd1 vssd1 vccd1 vccd1 hold2206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 _14799_/X vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08861_ _09015_/A hold305/X vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__and2_1
Xhold2228 _08063_/X vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2239 _15138_/X vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1505 _17907_/Q vssd1 vssd1 vccd1 vccd1 hold1505/X sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ _16286_/Q _07810_/Y hold2012/X _09339_/B vssd1 vssd1 vccd1 vccd1 _07812_/Y
+ sky130_fd_sc_hd__a31oi_1
Xhold1516 _08273_/X vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ _15482_/A hold666/X vssd1 vssd1 vccd1 vccd1 _16016_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1527 _17869_/Q vssd1 vssd1 vccd1 vccd1 hold1527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _15875_/Q vssd1 vssd1 vccd1 vccd1 hold1538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1549 _17826_/Q vssd1 vssd1 vccd1 vccd1 hold1549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09413_ _07804_/A _09456_/C _15264_/A _09412_/X vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09344_ _15217_/A hold469/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09363_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09275_ _15551_/A hold1311/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ hold1418/X _08209_/B _08225_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08157_ hold203/X hold690/X vssd1 vssd1 vccd1 vccd1 _08170_/S sky130_fd_sc_hd__nand2b_4
XFILLER_0_71_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ _14774_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4120 _10942_/X vssd1 vssd1 vccd1 vccd1 _16804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4131 _16582_/Q vssd1 vssd1 vccd1 vccd1 hold4131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4142 _13390_/X vssd1 vssd1 vccd1 vccd1 _17583_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4153 _17186_/Q vssd1 vssd1 vccd1 vccd1 hold4153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4164 _16608_/Q vssd1 vssd1 vccd1 vccd1 hold4164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4175 _16691_/Q vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3430 _17458_/Q vssd1 vssd1 vccd1 vccd1 hold3430/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _13246_/A _09954_/A _10049_/X vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4186 _13663_/X vssd1 vssd1 vccd1 vccd1 _17674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3441 _12241_/X vssd1 vssd1 vccd1 vccd1 _17237_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3452 _16357_/Q vssd1 vssd1 vccd1 vccd1 hold3452/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4197 _17716_/Q vssd1 vssd1 vccd1 vccd1 hold4197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3463 _13504_/X vssd1 vssd1 vccd1 vccd1 _17621_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3474 _17621_/Q vssd1 vssd1 vccd1 vccd1 hold3474/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3485 _13378_/X vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2740 _09157_/X vssd1 vssd1 vccd1 vccd1 _16191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2751 _14641_/X vssd1 vssd1 vccd1 vccd1 _18111_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3496 _17280_/Q vssd1 vssd1 vccd1 vccd1 hold3496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2762 _08220_/X vssd1 vssd1 vccd1 vccd1 _15746_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2773 _08222_/X vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2784 _16250_/Q vssd1 vssd1 vccd1 vccd1 hold2784/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2795 _17865_/Q vssd1 vssd1 vccd1 vccd1 hold2795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ _13761_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10952_ hold3010/X _16808_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13671_ _13698_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10883_ hold426/X _16785_/Q _11168_/C vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15410_ hold93/X _15486_/A2 _09357_/B _16070_/Q vssd1 vssd1 vccd1 vccd1 _15410_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ hold2061/X _17385_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__mux2_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _18389_/CLK _16390_/D vssd1 vssd1 vccd1 vccd1 _16390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ _09424_/B _15477_/A2 _15487_/B1 hold549/X _15340_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12553_ hold2622/X hold3593/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18060_ _18060_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11504_ hold1589/X _16992_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__mux2_1
X_15272_ _15480_/A _15272_/B _15272_/C _15272_/D vssd1 vssd1 vccd1 vccd1 _15272_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _17335_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ _17889_/CLK _17011_/D vssd1 vssd1 vccd1 vccd1 _17011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ hold1895/X _14216_/Y _14222_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _14223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ hold2854/X hold3910/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_230_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18123_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ hold1699/X _16946_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__mux2_1
X_14154_ _15553_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13105_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__and2_1
X_10317_ _10554_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11297_ hold697/X hold4689/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__mux2_1
X_14085_ hold2903/X _14094_/B _14084_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _14085_/X
+ sky130_fd_sc_hd__o211a_1
X_13036_ hold960/X _13035_/X hold957/A vssd1 vssd1 vccd1 vccd1 hold961/A sky130_fd_sc_hd__mux2_1
XFILLER_0_237_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10248_ _10536_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__or2_1
X_17913_ _18006_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _17876_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
X_10179_ _10563_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17775_ _17775_/CLK _17775_/D vssd1 vssd1 vccd1 vccd1 _17775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14987_ hold3191/X hold514/X _14986_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _14987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16726_ _18226_/CLK _16726_/D vssd1 vssd1 vccd1 vccd1 _16726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ _14726_/A hold2559/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16657_ _18213_/CLK _16657_/D vssd1 vssd1 vccd1 vccd1 _16657_/Q sky130_fd_sc_hd__dfxtp_1
X_13869_ hold3629/X _13773_/A _13868_/X vssd1 vssd1 vccd1 vccd1 _13869_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _18447_/CLK _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16588_ _18144_/CLK _16588_/D vssd1 vssd1 vccd1 vccd1 _16588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18327_ _18327_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15539_ _15539_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_389_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17171_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09060_ hold498/X hold541/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold542/A sky130_fd_sc_hd__mux2_1
X_18258_ _18360_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_318_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17970_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08011_ _15525_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17209_ _17273_/CLK _17209_/D vssd1 vssd1 vccd1 vccd1 _17209_/Q sky130_fd_sc_hd__dfxtp_1
X_18189_ _18221_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold602 hold602/A vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 hold613/A vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 hold624/A vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 hold635/A vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold646 hold646/A vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 hold657/A vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 hold668/A vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold679 hold679/A vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ hold964/X hold5090/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ _12424_/A hold711/X vssd1 vssd1 vccd1 vccd1 _16074_/D sky130_fd_sc_hd__and2_1
Xhold2003 _14827_/X vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09893_ hold2284/X hold3768/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__mux2_1
Xhold2014 _07825_/X vssd1 vssd1 vccd1 vccd1 _17751_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2025 _16166_/Q vssd1 vssd1 vccd1 vccd1 hold2025/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2036 _09161_/X vssd1 vssd1 vccd1 vccd1 _16193_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 hold1302/A vssd1 vssd1 vccd1 vccd1 _15203_/A sky130_fd_sc_hd__buf_12
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 _15796_/Q vssd1 vssd1 vccd1 vccd1 hold2047/X sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ hold353/X hold493/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__mux2_1
Xhold1313 _18307_/Q vssd1 vssd1 vccd1 vccd1 hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _17796_/Q vssd1 vssd1 vccd1 vccd1 hold2058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 _09407_/X vssd1 vssd1 vccd1 vccd1 _16289_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _14091_/X vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 hold1335/A vssd1 vssd1 vccd1 vccd1 _14974_/A sky130_fd_sc_hd__clkbuf_16
Xhold1346 _18080_/Q vssd1 vssd1 vccd1 vccd1 hold1346/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1357 _08423_/X vssd1 vssd1 vccd1 vccd1 hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ hold607/X _16008_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold608/A sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1368 _07858_/X vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1379 _15802_/Q vssd1 vssd1 vccd1 vccd1 hold1379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_178_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09327_ _15169_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ _12738_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _16240_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ _14878_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09189_ hold2063/X _09218_/B _09188_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _09189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ hold3850/X _11124_/A _11219_/X vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11151_ hold3262/X _11631_/A _11150_/X vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ hold4791/X _10598_/B _10101_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10102_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11082_/X sky130_fd_sc_hd__or2_1
XTAP_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3260 _12524_/X vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _10603_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _16501_/D sky130_fd_sc_hd__nor2_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ _14910_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__or2_1
Xhold3271 _17506_/Q vssd1 vssd1 vccd1 vccd1 hold3271/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3282 _17490_/Q vssd1 vssd1 vccd1 vccd1 hold3282/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15890_ _17344_/CLK _15890_/D vssd1 vssd1 vccd1 vccd1 hold625/A sky130_fd_sc_hd__dfxtp_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3293 _12614_/X vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2570 _18010_/Q vssd1 vssd1 vccd1 vccd1 hold2570/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ hold2778/X _14828_/B _14840_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2581 _18040_/Q vssd1 vssd1 vccd1 vccd1 hold2581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2592 _15673_/Q vssd1 vssd1 vccd1 vccd1 hold2592/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1880 _14508_/X vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17560_ _17725_/CLK _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
X_14772_ _15004_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14772_/Y sky130_fd_sc_hd__nand2_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1891 input67/X vssd1 vssd1 vccd1 vccd1 hold1891/X sky130_fd_sc_hd__dlygate4sd3_1
X_11984_ hold1485/X _17152_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16511_ _18294_/CLK _16511_/D vssd1 vssd1 vccd1 vccd1 _16511_/Q sky130_fd_sc_hd__dfxtp_1
X_13723_ hold5759/X _13829_/B _13722_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17491_ _17491_/CLK _17491_/D vssd1 vssd1 vccd1 vccd1 _17491_/Q sky130_fd_sc_hd__dfxtp_1
X_10935_ _11670_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16442_ _18327_/CLK _16442_/D vssd1 vssd1 vccd1 vccd1 _16442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ hold3509/X _13883_/B _13653_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _11136_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12605_ hold3561/X _12604_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12605_/X sky130_fd_sc_hd__mux2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _18356_/CLK _16373_/D vssd1 vssd1 vccd1 vccd1 _16373_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ hold4344/X _13856_/B _13584_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10797_ _11082_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18112_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15324_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__and2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12536_ hold3274/X _12535_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_411_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17769_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _18043_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ _15255_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__or2_1
X_12467_ hold98/X _12509_/A2 _12507_/A3 _12466_/X _09055_/A vssd1 vssd1 vccd1 vccd1
+ hold99/A sky130_fd_sc_hd__o311a_1
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ _14330_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11418_ _11706_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__or2_1
X_15186_ hold1387/X _15221_/B _15185_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _15186_/X
+ sky130_fd_sc_hd__o211a_1
X_12398_ _12438_/A _12398_/B vssd1 vssd1 vccd1 vccd1 _17292_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14137_ hold1610/X _14142_/B _14136_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14137_/X
+ sky130_fd_sc_hd__o211a_1
X_11349_ _11553_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14068_ _14246_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ hold952/X _13019_/B hold918/X hold930/X vssd1 vssd1 vccd1 vccd1 hold953/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _18062_/CLK _17827_/D vssd1 vssd1 vccd1 vccd1 _17827_/Q sky130_fd_sc_hd__dfxtp_1
X_08560_ hold118/X _15904_/Q _08592_/S vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__mux2_1
XFILLER_0_234_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17758_ _17886_/CLK _17758_/D vssd1 vssd1 vccd1 vccd1 _17758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16709_ _18070_/CLK _16709_/D vssd1 vssd1 vccd1 vccd1 _16709_/Q sky130_fd_sc_hd__dfxtp_1
X_08491_ hold2231/X _08486_/B _08490_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08491_/X
+ sky130_fd_sc_hd__o211a_1
X_17689_ _17689_/CLK _17689_/D vssd1 vssd1 vccd1 vccd1 _17689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09112_ _15553_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_152_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16095_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _12444_/A hold545/X vssd1 vssd1 vccd1 vccd1 _16138_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold410 hold410/A vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold432 hold432/A vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold443/A vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 hold74/X vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__buf_4
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 hold465/A vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 hold476/A vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 hold77/X vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__buf_4
Xfanout901 hold746/X vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__buf_12
X_09945_ _10191_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__or2_1
Xfanout912 _15173_/A vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout923 hold998/X vssd1 vssd1 vccd1 vccd1 hold999/A sky130_fd_sc_hd__buf_6
Xfanout934 hold1015/X vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__clkbuf_16
Xfanout945 hold1152/X vssd1 vssd1 vccd1 vccd1 hold1112/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _10470_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__or2_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 hold1149/X vssd1 vssd1 vccd1 vccd1 hold1150/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _16233_/Q vssd1 vssd1 vccd1 vccd1 hold1121/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _15672_/Q vssd1 vssd1 vccd1 vccd1 hold1132/X sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _12416_/A hold450/X vssd1 vssd1 vccd1 vccd1 _16032_/D sky130_fd_sc_hd__and2_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _15173_/X vssd1 vssd1 vccd1 vccd1 hold1143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 la_data_in[23] vssd1 vssd1 vccd1 vccd1 hold1154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1165 _08176_/X vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1176 _16151_/Q vssd1 vssd1 vccd1 vccd1 hold1176/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _08099_/X vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08758_ _15304_/A hold843/X vssd1 vssd1 vccd1 vccd1 _15999_/D sky130_fd_sc_hd__and2_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _13016_/X vssd1 vssd1 vccd1 vccd1 _17516_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ hold271/X hold326/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10720_ hold5148/X _11207_/B _10719_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _10720_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10651_ _18461_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _16707_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_180_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _11194_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _16684_/D sky130_fd_sc_hd__nor2_1
X_13370_ _15866_/Q hold3697/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_192_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ hold4719/X _13794_/A _12320_/X vssd1 vssd1 vccd1 vccd1 _12321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15040_ _15052_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _18303_/D sky130_fd_sc_hd__and2_1
X_12252_ _13773_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _16891_/D sky130_fd_sc_hd__nor2_1
X_12183_ _13461_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ hold4155/X _11156_/B _11133_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _11134_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16991_ _17869_/CLK _16991_/D vssd1 vssd1 vccd1 vccd1 _16991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15942_ _17332_/CLK _15942_/D vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__dfxtp_1
X_11065_ hold5368/X _11159_/B _11064_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _11065_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3090 _18114_/Q vssd1 vssd1 vccd1 vccd1 hold3090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ _16496_/Q _10034_/B _10034_/C vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__and3_1
XFILLER_0_200_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _17712_/CLK _15873_/D vssd1 vssd1 vccd1 vccd1 _15873_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _14878_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__nand2_1
X_17612_ _17612_/CLK _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17543_ _18390_/CLK _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ hold3143/X _14774_/B _14754_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14755_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11967_ _12231_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13706_ hold2214/X hold4149/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__mux2_1
X_10918_ hold4513/X _11210_/B _10917_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__o211a_1
X_17474_ _17478_/CLK _17474_/D vssd1 vssd1 vccd1 vccd1 _17474_/Q sky130_fd_sc_hd__dfxtp_1
X_14686_ _14794_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11898_ _13782_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16425_ _18366_/CLK _16425_/D vssd1 vssd1 vccd1 vccd1 _16425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13637_ hold2609/X _17666_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10849_ hold5487/X _11156_/B _10848_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16356_ _18375_/CLK _16356_/D vssd1 vssd1 vccd1 vccd1 _16356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13568_ hold1340/X hold4413/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15307_ hold637/X _15487_/A2 _15484_/B1 hold771/X _15306_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _12531_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _17349_/D sky130_fd_sc_hd__and2_1
X_16287_ _18460_/CLK _16287_/D vssd1 vssd1 vccd1 vccd1 _16287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13499_ hold2611/X _17620_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13500_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5409 _16816_/Q vssd1 vssd1 vccd1 vccd1 hold5409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ _18026_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ hold588/X _15484_/A2 _09392_/D hold704/X vssd1 vssd1 vccd1 vccd1 _15238_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4708 _11217_/Y vssd1 vssd1 vccd1 vccd1 _11218_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4719 _17104_/Q vssd1 vssd1 vccd1 vccd1 hold4719/X sky130_fd_sc_hd__dlygate4sd3_1
X_15169_ _15169_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15169_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout208 fanout246/X vssd1 vssd1 vccd1 vccd1 _12052_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_26_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout219 _10019_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__clkbuf_8
X_07991_ hold1691/X _07991_/A2 _07990_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _07991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09730_ hold4501/X _11201_/B _09729_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _09730_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09661_ hold4705/X _10055_/B _09660_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09661_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ _09053_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _15928_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ hold5162/X _10468_/A2 _09591_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09592_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08543_ _09063_/A hold155/X vssd1 vssd1 vccd1 vccd1 _15895_/D sky130_fd_sc_hd__and2_1
XFILLER_0_194_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_333_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17274_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08474_ _15207_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ hold454/X hold674/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__mux2_1
Xhold5910 _16319_/Q vssd1 vssd1 vccd1 vccd1 hold5910/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5921 _17535_/Q vssd1 vssd1 vccd1 vccd1 hold5921/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5932 _17532_/Q vssd1 vssd1 vccd1 vccd1 hold5932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5943 _17531_/Q vssd1 vssd1 vccd1 vccd1 hold5943/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5954 data_in[9] vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5965 hold6029/X vssd1 vssd1 vccd1 vccd1 hold5965/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__clkbuf_16
Xhold251 input30/X vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5976 _18367_/Q vssd1 vssd1 vccd1 vccd1 hold5976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold262 input20/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__buf_1
XFILLER_0_229_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5987 _18368_/Q vssd1 vssd1 vccd1 vccd1 hold5987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold273 hold364/X vssd1 vssd1 vccd1 vccd1 hold365/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5998 _18273_/Q vssd1 vssd1 vccd1 vccd1 hold5998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout720 _14434_/C1 vssd1 vssd1 vccd1 vccd1 _14366_/A sky130_fd_sc_hd__buf_4
Xfanout731 _12424_/A vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__buf_4
Xfanout742 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__buf_4
X_09928_ hold5527/X _11201_/B _09927_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09928_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout753 fanout770/X vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__buf_4
Xfanout764 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__buf_4
Xfanout775 _08125_/A vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__buf_4
Xfanout786 _14348_/A vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__buf_4
X_09859_ hold3655/X _10565_/B _09858_/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 _09859_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout797 _15056_/A vssd1 vssd1 vccd1 vccd1 _15194_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_213_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12870_ _12870_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _17466_/D sky130_fd_sc_hd__and2_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11821_ hold5290/X _12299_/B _11820_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ hold2840/X _14541_/B _14539_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14540_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _12340_/A _11752_/B vssd1 vssd1 vccd1 vccd1 _17074_/D sky130_fd_sc_hd__nor2_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ hold3082/X hold4678/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14471_ _14758_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14471_/X sky130_fd_sc_hd__or2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ hold5034/X _12317_/B _11682_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11683_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16210_ _17446_/CLK _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13422_ _13713_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10634_ _16702_/Q _11180_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _10634_/X sky130_fd_sc_hd__and3_1
X_17190_ _17623_/CLK _17190_/D vssd1 vssd1 vccd1 vccd1 _17190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16141_ _17340_/CLK _16141_/D vssd1 vssd1 vccd1 vccd1 _16141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13353_ _13698_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__or2_1
X_10565_ _16679_/Q _10565_/B _10565_/C vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__and3_1
XFILLER_0_88_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12304_ _13825_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _17258_/D sky130_fd_sc_hd__nor2_1
X_16072_ _17303_/CLK _16072_/D vssd1 vssd1 vccd1 vccd1 hold848/A sky130_fd_sc_hd__dfxtp_1
X_13284_ hold4707/X _13283_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10496_ hold2989/X hold3326/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15023_ _15131_/A hold1072/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15023_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12235_ hold5328/X _12329_/B _12234_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _12235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ hold5427/X _13862_/B _12165_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12166_/X
+ sky130_fd_sc_hd__o211a_1
X_11117_ hold2840/X _16863_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12097_ hold5383/X _12293_/B _12096_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16974_ _17852_/CLK _16974_/D vssd1 vssd1 vccd1 vccd1 _16974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _17314_/CLK _15925_/D vssd1 vssd1 vccd1 vccd1 hold628/A sky130_fd_sc_hd__dfxtp_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ hold797/X hold4346/X _11147_/C vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _17677_/CLK _15856_/D vssd1 vssd1 vccd1 vccd1 _15856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14807_ hold3053/X _14828_/B _14806_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14807_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15787_ _17726_/CLK _15787_/D vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ _12999_/A _12999_/B vssd1 vssd1 vccd1 vccd1 _17509_/D sky130_fd_sc_hd__and2_1
XFILLER_0_231_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17526_ _17534_/CLK _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_1
X_14738_ _15131_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ _18432_/CLK _17457_/D vssd1 vssd1 vccd1 vccd1 _17457_/Q sky130_fd_sc_hd__dfxtp_1
X_14669_ hold2532/X _14664_/B _14668_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16408_ _18319_/CLK _16408_/D vssd1 vssd1 vccd1 vccd1 _16408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08190_ hold1130/X _08213_/B _08189_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17388_ _18453_/CLK _17388_/D vssd1 vssd1 vccd1 vccd1 _17388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ _18316_/CLK _16339_/D vssd1 vssd1 vccd1 vccd1 _16339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5206 _16512_/Q vssd1 vssd1 vccd1 vccd1 hold5206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5217 _11530_/X vssd1 vssd1 vccd1 vccd1 _17000_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5228 _17031_/Q vssd1 vssd1 vccd1 vccd1 hold5228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5239 _13699_/X vssd1 vssd1 vccd1 vccd1 _17686_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4505 _17681_/Q vssd1 vssd1 vccd1 vccd1 hold4505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18009_ _18041_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4516 _11704_/X vssd1 vssd1 vccd1 vccd1 _17058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4527 hold5889/X vssd1 vssd1 vccd1 vccd1 hold5890/A sky130_fd_sc_hd__buf_6
XFILLER_0_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4538 _11125_/X vssd1 vssd1 vccd1 vccd1 _16865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3804 _16847_/Q vssd1 vssd1 vccd1 vccd1 hold3804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4549 _17058_/Q vssd1 vssd1 vccd1 vccd1 hold4549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3815 _17431_/Q vssd1 vssd1 vccd1 vccd1 hold3815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3826 _12345_/Y vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3837 _17191_/Q vssd1 vssd1 vccd1 vccd1 hold3837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3848 _17629_/Q vssd1 vssd1 vccd1 vccd1 hold3848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3859 _09745_/X vssd1 vssd1 vccd1 vccd1 _16405_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07974_ _15543_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09713_ hold2898/X hold3970/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09644_ hold1398/X _16372_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09575_ hold1981/X _13262_/A _10055_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__mux2_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ hold312/X hold725/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold726/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08457_ hold2643/X _08488_/B _08456_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08457_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _14443_/A hold1260/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _10524_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ _12430_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _16121_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5740 _13450_/X vssd1 vssd1 vccd1 vccd1 _17603_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10281_ _10560_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__or2_1
Xhold5751 _17728_/Q vssd1 vssd1 vccd1 vccd1 hold5751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5762 _13441_/X vssd1 vssd1 vccd1 vccd1 _17600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5773 hold5927/X vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5784 hold5784/A vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ hold1285/X hold5100/X _13412_/S vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__mux2_1
Xhold5795 hold5918/X vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout550 _08283_/Y vssd1 vssd1 vccd1 vccd1 _08336_/A2 sky130_fd_sc_hd__buf_8
Xfanout561 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout572 _07829_/Y vssd1 vssd1 vccd1 vccd1 _07865_/B sky130_fd_sc_hd__buf_8
Xfanout583 _13053_/X vssd1 vssd1 vccd1 vccd1 _13302_/B sky130_fd_sc_hd__buf_6
X_13971_ hold2369/X _13995_/A2 _13970_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _13971_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout594 _12826_/S vssd1 vssd1 vccd1 vccd1 _12913_/S sky130_fd_sc_hd__buf_6
X_15710_ _17278_/CLK hold369/X vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_255_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18230_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12922_ hold1714/X hold3290/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux2_1
X_16690_ _18214_/CLK _16690_/D vssd1 vssd1 vccd1 vccd1 _16690_/Q sky130_fd_sc_hd__dfxtp_1
X_15641_ _17153_/CLK _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ hold2757/X _17462_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18360_ _18360_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11804_ hold1163/X _17092_/Q _12029_/S vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__mux2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _17274_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12784_ hold1050/X _17439_/Q _12808_/S vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__mux2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17311_ _17335_/CLK _17311_/D vssd1 vssd1 vccd1 vccd1 _17311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14988_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__or2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18291_ _18387_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _17069_/Q _11738_/B _11738_/C vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17274_/CLK _17242_/D vssd1 vssd1 vccd1 vccd1 _17242_/Q sky130_fd_sc_hd__dfxtp_1
X_14454_ hold1901/X _14482_/A2 _14453_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ hold2683/X _17046_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13405_ hold4313/X _13883_/B _13404_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13405_/X
+ sky130_fd_sc_hd__o211a_1
X_10617_ hold4655/X _11103_/A _10616_/X vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__a21oi_1
X_17173_ _17269_/CLK _17173_/D vssd1 vssd1 vccd1 vccd1 _17173_/Q sky130_fd_sc_hd__dfxtp_1
X_14385_ _14726_/A hold2664/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ hold1527/X hold4277/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _17347_/CLK _16124_/D vssd1 vssd1 vccd1 vccd1 _16124_/Q sky130_fd_sc_hd__dfxtp_1
X_13336_ hold4081/X _13814_/B _13335_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _13336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10998_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16055_ _16089_/CLK _16055_/D vssd1 vssd1 vccd1 vccd1 hold473/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13267_ _13266_/X _16926_/Q _13267_/S vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__mux2_1
X_10479_ _11082_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__or2_1
X_15006_ _15221_/A hold514/X vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nand2_1
X_12218_ hold1444/X _17230_/Q _12314_/C vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__mux2_1
X_13198_ _13198_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12149_ hold2162/X _17207_/Q _12365_/C vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1709 _14067_/X vssd1 vssd1 vccd1 vccd1 _17836_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16957_ _17890_/CLK _16957_/D vssd1 vssd1 vccd1 vccd1 _16957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15908_ _17326_/CLK _15908_/D vssd1 vssd1 vccd1 vccd1 hold651/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16888_ _18226_/CLK _16888_/D vssd1 vssd1 vccd1 vccd1 _16888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15839_ _17666_/CLK _15839_/D vssd1 vssd1 vccd1 vccd1 _15839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09360_ _09366_/A _09360_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09362_/C sky130_fd_sc_hd__nor3_4
XFILLER_0_34_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _15535_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _17509_/CLK _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09291_ _14972_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _14246_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08242_/X sky130_fd_sc_hd__or2_1
XANTENNA_24 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 _14862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_46 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_57 hold607/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18305_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08173_ hold203/X _15182_/A vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_68 hold998/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_79 hold5866/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5003 _11710_/X vssd1 vssd1 vccd1 vccd1 _17060_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5014 _16935_/Q vssd1 vssd1 vccd1 vccd1 hold5014/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5025 _11830_/X vssd1 vssd1 vccd1 vccd1 _17100_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5036 _17060_/Q vssd1 vssd1 vccd1 vccd1 hold5036/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4302 _12079_/X vssd1 vssd1 vccd1 vccd1 _17183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5047 _10693_/X vssd1 vssd1 vccd1 vccd1 _16721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5058 _16703_/Q vssd1 vssd1 vccd1 vccd1 hold5058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4313 _17620_/Q vssd1 vssd1 vccd1 vccd1 hold4313/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput120 hold5876/X vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_12
Xoutput131 hold5866/X vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_12
Xhold4324 _13462_/X vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5069 _11766_/Y vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__dlygate4sd3_1
Xoutput142 _13029_/A vssd1 vssd1 vccd1 vccd1 load_status[2] sky130_fd_sc_hd__buf_12
XFILLER_0_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4335 _13402_/X vssd1 vssd1 vccd1 vccd1 _17587_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4346 _16840_/Q vssd1 vssd1 vccd1 vccd1 hold4346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3601 _11730_/Y vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3612 _12333_/Y vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4357 _13372_/X vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3623 _17118_/Q vssd1 vssd1 vccd1 vccd1 hold3623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4368 _17088_/Q vssd1 vssd1 vccd1 vccd1 hold4368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3634 _13815_/Y vssd1 vssd1 vccd1 vccd1 _13816_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4379 _11605_/X vssd1 vssd1 vccd1 vccd1 _17025_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3645 _17106_/Q vssd1 vssd1 vccd1 vccd1 hold3645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2900 _14339_/X vssd1 vssd1 vccd1 vccd1 _17967_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3656 _09859_/X vssd1 vssd1 vccd1 vccd1 _16443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2911 _17886_/Q vssd1 vssd1 vccd1 vccd1 hold2911/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2922 _14309_/X vssd1 vssd1 vccd1 vccd1 _17952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3667 _13839_/Y vssd1 vssd1 vccd1 vccd1 _13840_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3678 _10147_/X vssd1 vssd1 vccd1 vccd1 _16539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2933 _16269_/Q vssd1 vssd1 vccd1 vccd1 hold2933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3689 _16555_/Q vssd1 vssd1 vccd1 vccd1 hold3689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 _14550_/X vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2955 _18094_/Q vssd1 vssd1 vccd1 vccd1 hold2955/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2966 _17978_/Q vssd1 vssd1 vccd1 vccd1 hold2966/X sky130_fd_sc_hd__dlygate4sd3_1
X_07957_ hold3102/X _07991_/A2 _07956_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2977 _08071_/X vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2988 _08012_/X vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2999 _15810_/Q vssd1 vssd1 vccd1 vccd1 hold2999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07888_ hold915/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07888_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09627_ _09963_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ _09960_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09558_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08509_ _15513_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _13048_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _11712_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11643_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ hold3326/X _10628_/B _10401_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _10402_/X
+ sky130_fd_sc_hd__o211a_1
X_14170_ _15515_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14170_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ _11670_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13121_ _13121_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__and2_1
XFILLER_0_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ hold5330/X _10619_/B _10332_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5570 _11290_/X vssd1 vssd1 vccd1 vccd1 _16920_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13052_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13052_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_0_237_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10264_ hold4169/X _10628_/B _10263_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10264_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5581 _16979_/Q vssd1 vssd1 vccd1 vccd1 hold5581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5592 _10762_/X vssd1 vssd1 vccd1 vccd1 _16744_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _13797_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or2_1
Xhold4880 _10195_/X vssd1 vssd1 vccd1 vccd1 _16555_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10195_ hold4879/X _10601_/B _10194_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10195_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4891 _16687_/Q vssd1 vssd1 vccd1 vccd1 hold4891/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_436_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17860_ _17860_/CLK _17860_/D vssd1 vssd1 vccd1 vccd1 _17860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16811_ _18012_/CLK _16811_/D vssd1 vssd1 vccd1 vccd1 _16811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ _17855_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout380 _14830_/B vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__buf_6
XFILLER_0_22_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout391 _14626_/Y vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13954_ _15515_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13954_/X sky130_fd_sc_hd__or2_1
X_16742_ _18039_/CLK _16742_/D vssd1 vssd1 vccd1 vccd1 _16742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12905_ hold3161/X _12904_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__mux2_1
X_16673_ _18229_/CLK _16673_/D vssd1 vssd1 vccd1 vccd1 _16673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13885_ _13888_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _17748_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18412_ _18413_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ _17179_/CLK _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ hold3355/X _12835_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__mux2_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _18363_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
X_15555_ _15555_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__or2_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12767_ hold4237/X _12766_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__mux2_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14506_ hold1416/X _14535_/B _14505_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14506_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _18380_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ hold4683/X _12204_/A _11717_/X vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__a21oi_1
X_15486_ hold308/X _15486_/A2 _09362_/C hold91/X vssd1 vssd1 vccd1 vccd1 _15486_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ hold3760/X _12697_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14437_ _15551_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__or2_1
X_17225_ _17257_/CLK _17225_/D vssd1 vssd1 vccd1 vccd1 _17225_/Q sky130_fd_sc_hd__dfxtp_1
Xinput11 input11/A vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_6
XFILLER_0_128_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11649_ _11652_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11649_/X sky130_fd_sc_hd__or2_1
Xinput22 input22/A vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_6
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput33 input33/A vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 input44/A vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17156_ _17188_/CLK _17156_/D vssd1 vssd1 vccd1 vccd1 _17156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14368_ _14368_/A _14368_/B vssd1 vssd1 vccd1 vccd1 _17981_/D sky130_fd_sc_hd__and2_1
Xinput55 input55/A vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold806 hold806/A vssd1 vssd1 vccd1 vccd1 input54/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _17330_/CLK _16107_/D vssd1 vssd1 vccd1 vccd1 hold656/A sky130_fd_sc_hd__dfxtp_1
Xhold817 hold817/A vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold828 hold828/A vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ hold2475/X hold4114/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold839 hold839/A vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ _17891_/CLK _17087_/D vssd1 vssd1 vccd1 vccd1 _17087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ hold5978/X hold756/X _14298_/X _14356_/A vssd1 vssd1 vccd1 vccd1 hold757/A
+ sky130_fd_sc_hd__o211a_1
X_16038_ _18408_/CLK _16038_/D vssd1 vssd1 vccd1 vccd1 hold827/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ hold140/X hold304/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_177_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18381_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2207 _09296_/X vssd1 vssd1 vccd1 vccd1 _16258_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2218 _17903_/Q vssd1 vssd1 vccd1 vccd1 hold2218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2229 _15740_/Q vssd1 vssd1 vccd1 vccd1 hold2229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07811_ hold952/X hold930/X hold918/X _13019_/B vssd1 vssd1 vccd1 vccd1 _07811_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1506 _14213_/X vssd1 vssd1 vccd1 vccd1 _17907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17293_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1517 _16253_/Q vssd1 vssd1 vccd1 vccd1 hold1517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08791_ hold498/X hold665/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold666/A sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17989_ _18052_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1528 _14135_/X vssd1 vssd1 vccd1 vccd1 _17869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _08493_/X vssd1 vssd1 vccd1 vccd1 _15875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ _09438_/B _16292_/Q vssd1 vssd1 vccd1 vccd1 _09412_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ _15559_/A _15231_/A hold531/A hold391/A vssd1 vssd1 vccd1 vccd1 _09352_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _12759_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _16248_/D sky130_fd_sc_hd__and2_1
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _15559_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08156_ hold752/A hold689/X hold764/X hold732/X vssd1 vssd1 vccd1 vccd1 hold690/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_16_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08087_ hold1917/X _08088_/B _08086_/Y _08145_/A vssd1 vssd1 vccd1 vccd1 _08087_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4110 _17242_/Q vssd1 vssd1 vccd1 vccd1 hold4110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4121 _17278_/Q vssd1 vssd1 vccd1 vccd1 hold4121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4132 _10180_/X vssd1 vssd1 vccd1 vccd1 _16550_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4143 _17218_/Q vssd1 vssd1 vccd1 vccd1 hold4143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4154 _11992_/X vssd1 vssd1 vccd1 vccd1 _17154_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4165 _10258_/X vssd1 vssd1 vccd1 vccd1 _16576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3420 _12848_/X vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3431 _17383_/Q vssd1 vssd1 vccd1 vccd1 hold3431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4176 _10507_/X vssd1 vssd1 vccd1 vccd1 _16659_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4187 _17236_/Q vssd1 vssd1 vccd1 vccd1 hold4187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3442 _17237_/Q vssd1 vssd1 vccd1 vccd1 hold3442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3453 _09505_/X vssd1 vssd1 vccd1 vccd1 _16325_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4198 _13693_/X vssd1 vssd1 vccd1 vccd1 _17684_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3464 _17201_/Q vssd1 vssd1 vccd1 vccd1 hold3464/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3475 _13408_/X vssd1 vssd1 vccd1 vccd1 _17589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2730 _07838_/X vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 _15687_/Q vssd1 vssd1 vccd1 vccd1 hold2741/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3486 _17016_/Q vssd1 vssd1 vccd1 vccd1 hold3486/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ hold145/X hold196/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__mux2_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2752 _16251_/Q vssd1 vssd1 vccd1 vccd1 hold2752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3497 _12274_/X vssd1 vssd1 vccd1 vccd1 _17248_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2763 _17854_/Q vssd1 vssd1 vccd1 vccd1 hold2763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2774 _18127_/Q vssd1 vssd1 vccd1 vccd1 hold2774/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2785 _15649_/Q vssd1 vssd1 vccd1 vccd1 hold2785/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2796 _14127_/X vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10951_ hold4457/X _11147_/B _10950_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10951_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13670_ hold3017/X _17677_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10882_ hold5409/X _11732_/B _10881_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _10882_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12870_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _17383_/D sky130_fd_sc_hd__and2_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ hold828/X _15486_/A2 _09357_/B hold847/X vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ _13002_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _17360_/D sky130_fd_sc_hd__and2_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11503_ hold4277/X _12344_/B _11502_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11503_/X
+ sky130_fd_sc_hd__o211a_1
X_15271_ _16291_/Q _15477_/A2 _15487_/B1 hold464/X _15270_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ hold83/X _12509_/A2 _12507_/A3 _12482_/X _15491_/A vssd1 vssd1 vccd1 vccd1
+ hold84/A sky130_fd_sc_hd__o311a_1
XFILLER_0_227_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17010_ _17888_/CLK _17010_/D vssd1 vssd1 vccd1 vccd1 _17010_/Q sky130_fd_sc_hd__dfxtp_1
X_14222_ _14972_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11434_ hold5062/X _12299_/B _11433_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ hold1483/X _14148_/B _14152_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11365_ hold4487/X _12338_/B _11364_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11365_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18436_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13104_ _13097_/X _13103_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17531_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_225_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10316_ hold1569/X _16596_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__mux2_1
X_14084_ _15537_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11296_ hold5519/X _12338_/B _11295_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13035_ _17523_/Q _13034_/X _13048_/A _13035_/D vssd1 vssd1 vccd1 vccd1 _13035_/X
+ sky130_fd_sc_hd__and4bb_1
X_17912_ _18006_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_1
X_10247_ hold1509/X hold4921/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_270_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18220_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17843_ _17975_/CLK _17843_/D vssd1 vssd1 vccd1 vccd1 _17843_/Q sky130_fd_sc_hd__dfxtp_1
X_10178_ hold1789/X _16550_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17774_ _17870_/CLK _17774_/D vssd1 vssd1 vccd1 vccd1 _17774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14986_ _15201_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _18054_/CLK _16725_/D vssd1 vssd1 vccd1 vccd1 _16725_/Q sky130_fd_sc_hd__dfxtp_1
X_13937_ _13943_/A _13937_/B vssd1 vssd1 vccd1 vccd1 _17774_/D sky130_fd_sc_hd__and2_1
XFILLER_0_187_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16656_ _18176_/CLK _16656_/D vssd1 vssd1 vccd1 vccd1 _16656_/Q sky130_fd_sc_hd__dfxtp_1
X_13868_ _17743_/Q _13868_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ _17444_/CLK _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_1
X_12819_ _12894_/A _12819_/B vssd1 vssd1 vccd1 vccd1 _17449_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16587_ _18175_/CLK _16587_/D vssd1 vssd1 vccd1 vccd1 _16587_/Q sky130_fd_sc_hd__dfxtp_1
X_13799_ hold1418/X hold3704/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18326_ _18382_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ hold2844/X _15547_/B _15537_/X _12657_/A vssd1 vssd1 vccd1 vccd1 _15538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15469_ _17322_/Q _09357_/A _09392_/B hold165/X _15468_/X vssd1 vssd1 vccd1 vccd1
+ _15471_/C sky130_fd_sc_hd__a221o_1
X_18257_ _18360_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08010_ hold1199/X _08029_/B _08009_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08010_/X
+ sky130_fd_sc_hd__o211a_1
X_17208_ _17274_/CLK _17208_/D vssd1 vssd1 vccd1 vccd1 _17208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18188_ _18220_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
Xhold603 hold603/A vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold614 hold614/A vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_358_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17639_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17139_ _17171_/CLK _17139_/D vssd1 vssd1 vccd1 vccd1 _17139_/Q sky130_fd_sc_hd__dfxtp_1
Xhold625 hold625/A vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 hold636/A vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 hold647/A vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold658 hold658/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ hold4797/X _10055_/B _09960_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09961_/X
+ sky130_fd_sc_hd__o211a_1
Xhold669 hold669/A vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ hold228/X hold710/X _08912_/S vssd1 vssd1 vccd1 vccd1 hold711/A sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09892_ hold5118/X _10034_/B _09891_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09892_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _15793_/Q vssd1 vssd1 vccd1 vccd1 hold2004/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 _15630_/Q vssd1 vssd1 vccd1 vccd1 hold2015/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2026 _09103_/X vssd1 vssd1 vccd1 vccd1 _16166_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08843_ _15324_/A hold673/X vssd1 vssd1 vccd1 vccd1 _16040_/D sky130_fd_sc_hd__and2_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _15808_/Q vssd1 vssd1 vccd1 vccd1 hold2037/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1303 _08250_/X vssd1 vssd1 vccd1 vccd1 hold1303/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2048 _08326_/X vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _15670_/Q vssd1 vssd1 vccd1 vccd1 hold1314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 _13983_/X vssd1 vssd1 vccd1 vccd1 _17796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 _16259_/Q vssd1 vssd1 vccd1 vccd1 hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1336 _14904_/X vssd1 vssd1 vccd1 vccd1 hold1336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _15394_/A hold423/X vssd1 vssd1 vccd1 vccd1 _16007_/D sky130_fd_sc_hd__and2_1
Xhold1347 _14577_/X vssd1 vssd1 vccd1 vccd1 _18080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 _08424_/X vssd1 vssd1 vccd1 vccd1 _15842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1369 _15637_/Q vssd1 vssd1 vccd1 vccd1 hold1369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18042_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09326_ hold2457/X _09338_/A2 _09325_/Y _12600_/A vssd1 vssd1 vccd1 vccd1 _09326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09257_ _15533_/A hold2662/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08208_ hold2229/X _08213_/B _08207_/Y _08143_/A vssd1 vssd1 vccd1 vccd1 _08208_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09188_ _15517_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08139_ _08139_/A hold241/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__and2_1
XFILLER_0_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11150_ _16874_/Q _11150_/B _11150_/C vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__and3_1
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10101_ _10563_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2_1
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ hold2577/X hold4703/X _11177_/C vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__mux2_1
XTAP_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3250 _17349_/Q vssd1 vssd1 vccd1 vccd1 hold3250/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _13198_/A _09960_/A _10031_/X vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__a21oi_1
Xhold3261 _17352_/Q vssd1 vssd1 vccd1 vccd1 hold3261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3272 _12989_/X vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3283 _17496_/Q vssd1 vssd1 vccd1 vccd1 hold3283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3294 _17484_/Q vssd1 vssd1 vccd1 vccd1 hold3294/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2560 _15583_/Q vssd1 vssd1 vccd1 vccd1 hold2560/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _15233_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__or2_1
Xhold2571 _14428_/X vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 _14490_/X vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2593 _08067_/X vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1870 _14225_/X vssd1 vssd1 vccd1 vccd1 _17912_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ hold2176/X _14774_/B _14770_/Y _14384_/A vssd1 vssd1 vccd1 vccd1 _14771_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1881 _16227_/Q vssd1 vssd1 vccd1 vccd1 hold1881/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11983_ hold4477/X _12344_/B _11982_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11983_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1892 _08467_/X vssd1 vssd1 vccd1 vccd1 _15862_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16510_ _18393_/CLK _16510_/D vssd1 vssd1 vccd1 vccd1 _16510_/Q sky130_fd_sc_hd__dfxtp_1
X_13722_ _13734_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13722_/X sky130_fd_sc_hd__or2_1
X_10934_ hold3124/X _16802_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_169_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17490_ _17491_/CLK _17490_/D vssd1 vssd1 vccd1 vccd1 _17490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16441_ _18384_/CLK _16441_/D vssd1 vssd1 vccd1 vccd1 _16441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _13788_/A _13653_/B vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10865_ hold2978/X hold3515/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ hold2876/X _17379_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__mux2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16372_ _18379_/CLK _16372_/D vssd1 vssd1 vccd1 vccd1 _16372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13584_ _13761_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ hold2753/X _16756_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _18143_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
X_15323_ _15490_/A1 _15315_/X _15322_/X _15490_/B1 hold5846/A vssd1 vssd1 vccd1 vccd1
+ _15323_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ hold1618/X hold3155/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15254_ _15414_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18042_ _18042_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12466_ _17326_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ hold2218/X _14202_/B _14204_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11417_ hold2153/X _16963_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__mux2_1
X_15185_ _15185_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_451_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17724_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12397_ hold174/X hold192/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _14529_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14136_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ hold1408/X hold5395/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14067_ hold1708/X _14107_/A2 _14066_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _14067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ hold1531/X hold5102/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ hold2535/X _13003_/Y _13017_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _17858_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _17887_/CLK _17757_/D vssd1 vssd1 vccd1 vccd1 _17757_/Q sky130_fd_sc_hd__dfxtp_1
X_14969_ hold1841/X _15004_/B _14968_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _14969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16708_ _18070_/CLK _16708_/D vssd1 vssd1 vccd1 vccd1 _16708_/Q sky130_fd_sc_hd__dfxtp_1
X_08490_ _14328_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17688_ _17726_/CLK _17688_/D vssd1 vssd1 vccd1 vccd1 _17688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16639_ _18123_/CLK _16639_/D vssd1 vssd1 vccd1 vccd1 _16639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ hold1252/X _09119_/A2 _09110_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09111_/X
+ sky130_fd_sc_hd__o211a_1
X_18309_ _18309_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09042_ hold228/X hold544/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold545/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold400 hold43/X vssd1 vssd1 vccd1 vccd1 input15/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_192_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18342_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold411 hold411/A vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold422 hold422/A vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold444 hold444/A vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold455 hold455/A vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold466 la_data_in[16] vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold477 hold477/A vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ hold1092/X hold5176/X _10190_/S vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__mux2_1
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 hold808/X vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__clkbuf_16
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _15173_/A vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout924 hold998/X vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout935 hold1015/X vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__buf_4
Xfanout946 hold1152/X vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__buf_8
X_09875_ hold1819/X hold3657/X _10565_/C vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _18436_/Q vssd1 vssd1 vccd1 vccd1 hold1100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 hold1151/X vssd1 vssd1 vccd1 vccd1 hold1152/A sky130_fd_sc_hd__buf_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ hold361/X hold449/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold450/A sky130_fd_sc_hd__mux2_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _09243_/X vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _08065_/X vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _15174_/X vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 hold1155/A vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 _16209_/Q vssd1 vssd1 vccd1 vccd1 hold1166/X sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ hold454/X hold842/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold843/A sky130_fd_sc_hd__mux2_1
Xhold1177 _09073_/X vssd1 vssd1 vccd1 vccd1 _16151_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1188 _15885_/Q vssd1 vssd1 vccd1 vccd1 hold1188/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1199 _15646_/Q vssd1 vssd1 vccd1 vccd1 hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08688_ _12531_/A hold650/X vssd1 vssd1 vccd1 vccd1 _15965_/D sky130_fd_sc_hd__and2_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ hold4617/X _10554_/A _10649_/X vssd1 vssd1 vccd1 vccd1 _10650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _15531_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10581_ hold4599/X _10563_/A _10580_/X vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _17264_/Q _12353_/B _13793_/S vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_209_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18143_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ hold2780/X hold3432/X _12251_/S vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11202_ hold4960/X _11106_/A _11201_/X vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12182_ hold2473/X hold4143/X _13556_/S vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__mux2_1
X_11133_ _11637_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16990_ _17867_/CLK _16990_/D vssd1 vssd1 vccd1 vccd1 _16990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15941_ _17301_/CLK _15941_/D vssd1 vssd1 vccd1 vccd1 hold539/A sky130_fd_sc_hd__dfxtp_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3080 _18004_/Q vssd1 vssd1 vccd1 vccd1 hold3080/X sky130_fd_sc_hd__dlygate4sd3_1
X_10015_ _11203_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _16495_/D sky130_fd_sc_hd__nor2_1
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3091 _14647_/X vssd1 vssd1 vccd1 vccd1 _18114_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _17711_/CLK _15872_/D vssd1 vssd1 vccd1 vccd1 _15872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 _08269_/X vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17611_ _17734_/CLK _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14823_ hold1579/X _14826_/B _14822_/Y _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14823_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17542_ _18318_/CLK _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14754_ _15201_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14754_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11966_ hold1241/X hold3436/X _12251_/S vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _11115_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__or2_1
X_13705_ hold3704/X _13814_/B _13704_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13705_/X
+ sky130_fd_sc_hd__o211a_1
X_14685_ hold1664/X _14720_/B _14684_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14685_/X
+ sky130_fd_sc_hd__o211a_1
X_17473_ _17877_/CLK _17473_/D vssd1 vssd1 vccd1 vccd1 _17473_/Q sky130_fd_sc_hd__dfxtp_1
X_11897_ hold1322/X hold3683/X _13877_/C vssd1 vssd1 vccd1 vccd1 _11898_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16424_ _18341_/CLK _16424_/D vssd1 vssd1 vccd1 vccd1 _16424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13636_ hold5717/X _13832_/B _13635_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13636_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_59_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_59_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_10848_ _11136_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16355_ _18266_/CLK _16355_/D vssd1 vssd1 vccd1 vccd1 _16355_/Q sky130_fd_sc_hd__dfxtp_1
X_13567_ hold4455/X _13883_/B _13566_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10779_ _11106_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ _17334_/Q _09362_/C _15485_/B1 hold436/X vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__a22o_1
X_12518_ hold3250/X _12517_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__mux2_1
X_16286_ _18237_/CLK _16286_/D vssd1 vssd1 vccd1 vccd1 _16286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13498_ hold4441/X _13880_/B _13497_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18025_ _18200_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ _16132_/Q _15487_/A2 _15484_/B1 _17307_/Q _15236_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/B sky130_fd_sc_hd__a221o_1
X_12449_ hold312/A _12509_/A2 _12507_/A3 _12448_/X _12424_/A vssd1 vssd1 vccd1 vccd1
+ hold102/A sky130_fd_sc_hd__o311a_1
XFILLER_0_48_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4709 _16447_/Q vssd1 vssd1 vccd1 vccd1 hold4709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15168_ hold2416/X _15167_/B _15167_/Y _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15168_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14119_ hold2274/X _14142_/B _14118_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15099_ _15099_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15099_/X sky130_fd_sc_hd__or2_1
Xfanout209 _10019_/B vssd1 vssd1 vccd1 vccd1 _11147_/B sky130_fd_sc_hd__buf_4
X_07990_ _14894_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09660_ _09960_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ hold47/X hold371/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__mux2_1
X_17809_ _17870_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09591_ _10467_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ hold17/X _15895_/Q _08592_/S vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08473_ hold2461/X _08486_/B _08472_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_373_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17680_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_302_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17767_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5900 _17521_/Q vssd1 vssd1 vccd1 vccd1 hold5900/X sky130_fd_sc_hd__dlygate4sd3_1
X_09025_ _12444_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _16129_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5911 _16906_/Q vssd1 vssd1 vccd1 vccd1 hold5911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5922 _17550_/Q vssd1 vssd1 vccd1 vccd1 hold5922/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5933 _17541_/Q vssd1 vssd1 vccd1 vccd1 hold5933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5944 _17555_/Q vssd1 vssd1 vccd1 vccd1 hold5944/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5955 data_in[22] vssd1 vssd1 vccd1 vccd1 hold604/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5966 data_in[23] vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5977 _15762_/Q vssd1 vssd1 vccd1 vccd1 hold5977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold62/X vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__clkbuf_8
Xhold5988 _18392_/Q vssd1 vssd1 vccd1 vccd1 hold5988/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5999 _15862_/Q vssd1 vssd1 vccd1 vccd1 hold5999/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold366/X vssd1 vssd1 vccd1 vccd1 hold367/A sky130_fd_sc_hd__buf_6
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout710 _13037_/A vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__buf_2
Xfanout721 _14434_/C1 vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout732 _12424_/A vssd1 vssd1 vccd1 vccd1 _12418_/A sky130_fd_sc_hd__clkbuf_4
X_09927_ _11106_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__or2_1
Xfanout743 _07787_/Y vssd1 vssd1 vccd1 vccd1 _14915_/C1 sky130_fd_sc_hd__buf_8
Xfanout754 fanout770/X vssd1 vssd1 vccd1 vccd1 _13657_/C1 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout765 _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__buf_4
XFILLER_0_226_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout776 fanout796/X vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__buf_4
X_09858_ _10470_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__or2_1
Xfanout787 _14348_/A vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__buf_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout798 _15056_/A vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__buf_4
XFILLER_0_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _09015_/A hold338/X vssd1 vssd1 vccd1 vccd1 _16023_/D sky130_fd_sc_hd__and2_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _11106_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__or2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _12204_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__or2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ hold4907/X _11658_/A _11750_/X vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ hold4825/X _11180_/B _10701_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10702_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ hold3031/X _14482_/A2 _14469_/X _14348_/A vssd1 vssd1 vccd1 vccd1 _14470_/X
+ sky130_fd_sc_hd__o211a_1
X_11682_ _12285_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ hold2699/X hold3942/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__mux2_1
X_10633_ _18461_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _16701_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16140_ _17315_/CLK _16140_/D vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13352_ hold2297/X hold5667/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ hold4329/X _10598_/B _10563_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _16678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12303_ hold3569/X _13716_/A _12302_/X vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__a21oi_1
X_16071_ _17320_/CLK _16071_/D vssd1 vssd1 vccd1 vccd1 hold740/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13283_ _13282_/X _16928_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10495_ hold4891/X _10649_/B _10494_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _15030_/A _15022_/B vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ _12261_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _11210_/A _11210_/B _11115_/X _14538_/C1 vssd1 vssd1 vccd1 vccd1 _11116_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12096_ _13797_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__or2_1
X_16973_ _17851_/CLK _16973_/D vssd1 vssd1 vccd1 vccd1 _16973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ _17299_/CLK _15924_/D vssd1 vssd1 vccd1 vccd1 hold759/A sky130_fd_sc_hd__dfxtp_1
X_11047_ hold4362/X _11147_/B _11046_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _11047_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 input9/A vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_6
XFILLER_0_204_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _17613_/CLK _15855_/D vssd1 vssd1 vccd1 vccd1 _15855_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14806_ _14984_/A _14830_/B vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15786_ _17650_/CLK _15786_/D vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ hold3276/X _12997_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__mux2_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _17525_/CLK _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14737_ hold1952/X _14772_/B _14736_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14737_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11949_ _13773_/A _11949_/B vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17456_ _18432_/CLK _17456_/D vssd1 vssd1 vccd1 vccd1 _17456_/Q sky130_fd_sc_hd__dfxtp_1
X_14668_ _15169_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ _18382_/CLK _16407_/D vssd1 vssd1 vccd1 vccd1 _16407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13619_ hold2004/X hold4073/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13620_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17387_ _18436_/CLK _17387_/D vssd1 vssd1 vccd1 vccd1 _17387_/Q sky130_fd_sc_hd__dfxtp_1
X_14599_ hold2884/X _14610_/B _14598_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16338_ _18351_/CLK _16338_/D vssd1 vssd1 vccd1 vccd1 _16338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5207 _09970_/X vssd1 vssd1 vccd1 vccd1 _16480_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16269_ _17370_/CLK _16269_/D vssd1 vssd1 vccd1 vccd1 _16269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5218 _17196_/Q vssd1 vssd1 vccd1 vccd1 hold5218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5229 _11527_/X vssd1 vssd1 vccd1 vccd1 _16999_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18040_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4506 _13588_/X vssd1 vssd1 vccd1 vccd1 _17649_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4517 _17217_/Q vssd1 vssd1 vccd1 vccd1 hold4517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4528 _15373_/X vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4539 _16833_/Q vssd1 vssd1 vccd1 vccd1 hold4539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3805 _10975_/X vssd1 vssd1 vccd1 vccd1 _16815_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3816 _12764_/X vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3827 _16467_/Q vssd1 vssd1 vccd1 vccd1 hold3827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3838 _12007_/X vssd1 vssd1 vccd1 vccd1 _17159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3849 _13432_/X vssd1 vssd1 vccd1 vccd1 _17597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07973_ hold2403/X _07978_/B _07972_/Y _15500_/A vssd1 vssd1 vccd1 vccd1 _07973_/X
+ sky130_fd_sc_hd__o211a_1
X_09712_ hold5362/X _11159_/B _09711_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _09712_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09643_ hold3359/X _10007_/B _09642_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09643_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09574_ hold5661/X _10070_/B _09573_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09574_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08525_ _15491_/A hold791/X vssd1 vssd1 vccd1 vccd1 _15887_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08456_ _14116_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08456_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _15825_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09008_ hold88/X hold92/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5730 _13738_/X vssd1 vssd1 vccd1 vccd1 _17699_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10280_ hold3067/X _16584_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__mux2_1
Xhold5741 _17665_/Q vssd1 vssd1 vccd1 vccd1 hold5741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5752 _13729_/X vssd1 vssd1 vccd1 vccd1 _17696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5763 hold5922/X vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5774 output89/X vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_12
Xhold5785 hold5932/X vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5796 output77/X vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout540 _08498_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__clkbuf_8
Xfanout551 _08260_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__buf_8
Xfanout562 _08043_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__buf_6
XFILLER_0_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout573 _07829_/Y vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__clkbuf_8
X_13970_ _15531_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__or2_1
Xfanout584 _13053_/X vssd1 vssd1 vccd1 vccd1 _13310_/B sky130_fd_sc_hd__buf_6
XFILLER_0_226_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout595 _12513_/X vssd1 vssd1 vccd1 vccd1 _12826_/S sky130_fd_sc_hd__clkbuf_4
X_12921_ _12921_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _17483_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _17215_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12921_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _17460_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _12367_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _17091_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_295_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18063_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12789_/A _12783_/B vssd1 vssd1 vccd1 vccd1 _17437_/D sky130_fd_sc_hd__and2_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _17777_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17330_/CLK _17310_/D vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__dfxtp_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ hold3213/X _14541_/B _14521_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14522_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11734_ _12310_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _17068_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_224_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18290_ _18322_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17241_ _17273_/CLK _17241_/D vssd1 vssd1 vccd1 vccd1 _17241_/Q sky130_fd_sc_hd__dfxtp_1
X_14453_ _14794_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__or2_1
X_11665_ hold5641/X _11789_/B _11664_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _11665_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ _10616_/A _11198_/B _11198_/C vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__and3_1
X_13404_ _13788_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__or2_1
X_14384_ _14384_/A _14384_/B vssd1 vssd1 vccd1 vccd1 _17989_/D sky130_fd_sc_hd__and2_1
X_17172_ _17236_/CLK _17172_/D vssd1 vssd1 vccd1 vccd1 _17172_/Q sky130_fd_sc_hd__dfxtp_1
X_11596_ hold4469/X _12338_/B _11595_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11596_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16123_ _16127_/CLK _16123_/D vssd1 vssd1 vccd1 vccd1 hold417/A sky130_fd_sc_hd__dfxtp_1
X_13335_ _13800_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ hold1001/X _16673_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _16077_/CLK _16054_/D vssd1 vssd1 vccd1 vccd1 hold419/A sky130_fd_sc_hd__dfxtp_1
X_13266_ _17584_/Q _17118_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13266_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10478_ hold1229/X _16650_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ hold1966/X _15004_/B _15004_/Y _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15005_/X
+ sky130_fd_sc_hd__o211a_1
X_12217_ hold5401/X _13862_/B _12216_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12217_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13197_ _13196_/X hold4637/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_202_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ hold5617/X _12338_/B _12147_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _12148_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12079_ hold4301/X _12374_/B _12078_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12079_/X
+ sky130_fd_sc_hd__o211a_1
X_16956_ _17834_/CLK _16956_/D vssd1 vssd1 vccd1 vccd1 _16956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15907_ _18423_/CLK _15907_/D vssd1 vssd1 vccd1 vccd1 hold694/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16887_ _18124_/CLK _16887_/D vssd1 vssd1 vccd1 vccd1 _16887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _17728_/CLK _15838_/D vssd1 vssd1 vccd1 vccd1 _15838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15769_ _17694_/CLK _15769_/D vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08310_ hold2836/X _08323_/B _08309_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _08310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17508_ _17508_/CLK _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_1
X_09290_ hold1327/X _09338_/A2 _09289_/X _12606_/A vssd1 vssd1 vccd1 vccd1 _09290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08241_ hold1706/X _08263_/A2 _08240_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08241_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_14 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _18434_/CLK _17439_/D vssd1 vssd1 vccd1 vccd1 _17439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_25 _14556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 _14862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_47 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 hold607/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ hold752/A hold689/A hold764/A hold732/A vssd1 vssd1 vccd1 vccd1 _15182_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_0_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_69 hold998/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5004 _16920_/Q vssd1 vssd1 vccd1 vccd1 hold5004/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5015 _11239_/X vssd1 vssd1 vccd1 vccd1 _16903_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5026 _16670_/Q vssd1 vssd1 vccd1 vccd1 hold5026/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18402_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5037 _11614_/X vssd1 vssd1 vccd1 vccd1 _17028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5048 _16422_/Q vssd1 vssd1 vccd1 vccd1 hold5048/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput110 hold5870/X vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4303 _17650_/Q vssd1 vssd1 vccd1 vccd1 hold4303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4314 _13405_/X vssd1 vssd1 vccd1 vccd1 _17588_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5059 _10543_/X vssd1 vssd1 vccd1 vccd1 _16671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput121 hold5885/X vssd1 vssd1 vccd1 vccd1 hold5886/A sky130_fd_sc_hd__buf_6
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput132 hold5842/X vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4325 _16961_/Q vssd1 vssd1 vccd1 vccd1 hold4325/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput143 hold5901/X vssd1 vssd1 vccd1 vccd1 load_status[3] sky130_fd_sc_hd__buf_12
Xhold4336 _16775_/Q vssd1 vssd1 vccd1 vccd1 hold4336/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17491_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4347 _10954_/X vssd1 vssd1 vccd1 vccd1 _16808_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3602 _17114_/Q vssd1 vssd1 vccd1 vccd1 hold3602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3613 _16415_/Q vssd1 vssd1 vccd1 vccd1 hold3613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4358 _17669_/Q vssd1 vssd1 vccd1 vccd1 hold4358/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3624 _12363_/Y vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4369 _11698_/X vssd1 vssd1 vccd1 vccd1 _17056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3635 _16411_/Q vssd1 vssd1 vccd1 vccd1 hold3635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2901 _16257_/Q vssd1 vssd1 vccd1 vccd1 hold2901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3646 _12327_/Y vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3657 _16449_/Q vssd1 vssd1 vccd1 vccd1 hold3657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2912 _14171_/X vssd1 vssd1 vccd1 vccd1 _17886_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3668 _16626_/Q vssd1 vssd1 vccd1 vccd1 hold3668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2923 _16190_/Q vssd1 vssd1 vccd1 vccd1 hold2923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2934 _09318_/X vssd1 vssd1 vccd1 vccd1 _16269_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3679 _16712_/Q vssd1 vssd1 vccd1 vccd1 hold3679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2945 _15734_/Q vssd1 vssd1 vccd1 vccd1 hold2945/X sky130_fd_sc_hd__dlygate4sd3_1
X_07956_ _15525_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_227_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2956 _14605_/X vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2967 _18219_/Q vssd1 vssd1 vccd1 vccd1 hold2967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2978 _17980_/Q vssd1 vssd1 vccd1 vccd1 hold2978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2989 _18212_/Q vssd1 vssd1 vccd1 vccd1 hold2989/X sky130_fd_sc_hd__dlygate4sd3_1
X_07887_ hold1269/X _07918_/B _07886_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _07887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09626_ hold3191/X hold3960/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09557_ hold1599/X _16343_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08508_ hold1088/X _08503_/Y _08507_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08508_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _17523_/Q _13035_/D vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08439_ _15553_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ hold2834/X _16974_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__mux2_1
X_10401_ _10497_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11381_ hold2711/X hold5623/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13113_/X _13119_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17533_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10332_ _10524_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13051_ _13051_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and2_1
Xhold5560 _10876_/X vssd1 vssd1 vccd1 vccd1 _16782_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10263_ _10527_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__or2_1
Xhold5571 _16370_/Q vssd1 vssd1 vccd1 vccd1 hold5571/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5582 _11371_/X vssd1 vssd1 vccd1 vccd1 _16947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5593 _16891_/Q vssd1 vssd1 vccd1 vccd1 hold5593/X sky130_fd_sc_hd__dlygate4sd3_1
X_12002_ hold1199/X hold5146/X _13412_/S vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4870 _10504_/X vssd1 vssd1 vccd1 vccd1 _16658_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10194_ _10488_/A _10194_/B vssd1 vssd1 vccd1 vccd1 _10194_/X sky130_fd_sc_hd__or2_1
Xhold4881 _16729_/Q vssd1 vssd1 vccd1 vccd1 hold4881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4892 _10495_/X vssd1 vssd1 vccd1 vccd1 _16655_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16810_ _18043_/CLK _16810_/D vssd1 vssd1 vccd1 vccd1 _16810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17790_ _17851_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout370 hold394/X vssd1 vssd1 vccd1 vccd1 _15069_/S sky130_fd_sc_hd__clkbuf_8
Xfanout381 _14788_/Y vssd1 vssd1 vccd1 vccd1 _14828_/B sky130_fd_sc_hd__buf_8
XFILLER_0_219_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _18070_/CLK _16741_/D vssd1 vssd1 vccd1 vccd1 _16741_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout392 _14543_/B vssd1 vssd1 vccd1 vccd1 _14553_/B sky130_fd_sc_hd__buf_6
XFILLER_0_199_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13953_ hold2888/X _13995_/A2 _13952_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _13953_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ hold2377/X _17479_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_236_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16672_ _18228_/CLK _16672_/D vssd1 vssd1 vccd1 vccd1 _16672_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_405_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17952_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13884_ hold3641/X _13788_/A _13883_/X vssd1 vssd1 vccd1 vccd1 _13884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18411_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15623_ _17153_/CLK _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ hold2808/X _17456_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18342_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ hold2632/X _15560_/A2 _15553_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _15554_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ hold1517/X hold3750/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ _15185_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__or2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18273_ _18273_/CLK hold515/X vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11717_ _17063_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__and3_1
X_15485_ hold90/X _15485_/A2 _15485_/B1 hold647/X vssd1 vssd1 vccd1 vccd1 _15485_/X
+ sky130_fd_sc_hd__a22o_1
X_12697_ hold2745/X _17410_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ _18447_/CLK _17224_/D vssd1 vssd1 vccd1 vccd1 _17224_/Q sky130_fd_sc_hd__dfxtp_1
X_14436_ hold2262/X _14433_/B _14435_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14436_/X
+ sky130_fd_sc_hd__o211a_1
X_11648_ hold2911/X _17040_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__mux2_1
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_6
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 input23/A vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_6
XFILLER_0_141_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput34 input34/A vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput45 input45/A vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_17155_ _17283_/CLK _17155_/D vssd1 vssd1 vccd1 vccd1 _17155_/Q sky130_fd_sc_hd__dfxtp_1
X_14367_ _15535_/A hold1903/X hold333/X vssd1 vssd1 vccd1 vccd1 _14368_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11579_ hold2240/X _17017_/Q _11594_/S vssd1 vssd1 vccd1 vccd1 _11580_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput56 input56/A vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_6
Xinput67 input67/A vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
Xhold807 input54/X vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16106_ _17329_/CLK _16106_/D vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold818 hold822/X vssd1 vssd1 vccd1 vccd1 hold823/A sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ hold5298/X _13798_/A2 _13317_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__o211a_1
Xhold829 hold829/A vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14298_ hold525/X _14336_/B vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__or2_1
X_17086_ _17900_/CLK _17086_/D vssd1 vssd1 vccd1 vccd1 _17086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _17293_/CLK _16037_/D vssd1 vssd1 vccd1 vccd1 hold387/A sky130_fd_sc_hd__dfxtp_1
X_13249_ _13249_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2208 _18324_/Q vssd1 vssd1 vccd1 vccd1 hold2208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2219 _14205_/X vssd1 vssd1 vccd1 vccd1 _17903_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07810_ _12412_/A _17751_/Q vssd1 vssd1 vccd1 vccd1 _07810_/Y sky130_fd_sc_hd__nand2_1
X_08790_ _15482_/A hold293/X vssd1 vssd1 vccd1 vccd1 _16015_/D sky130_fd_sc_hd__and2_1
Xhold1507 _17760_/Q vssd1 vssd1 vccd1 vccd1 hold1507/X sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ _18319_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1518 _09283_/X vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _18155_/Q vssd1 vssd1 vccd1 vccd1 hold1529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16939_ _18425_/CLK _16939_/D vssd1 vssd1 vccd1 vccd1 _16939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_146_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18366_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09411_ _07804_/A _09447_/A _15304_/A _09410_/X vssd1 vssd1 vccd1 vccd1 _09411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09273_ _15549_/A hold2178/X _09273_/S vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ hold1434/X _08209_/B _08223_/X _12747_/A vssd1 vssd1 vccd1 vccd1 _08224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _15004_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08086_/Y sky130_fd_sc_hd__nand2_1
Xhold4100 _10471_/X vssd1 vssd1 vccd1 vccd1 _16647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4111 _12160_/X vssd1 vssd1 vccd1 vccd1 _17210_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4122 _12268_/X vssd1 vssd1 vccd1 vccd1 _17246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4133 _17592_/Q vssd1 vssd1 vccd1 vccd1 hold4133/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4144 _12088_/X vssd1 vssd1 vccd1 vccd1 _17186_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4155 _16708_/Q vssd1 vssd1 vccd1 vccd1 hold4155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3410 _17415_/Q vssd1 vssd1 vccd1 vccd1 hold3410/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4166 _17658_/Q vssd1 vssd1 vccd1 vccd1 hold4166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3421 _17460_/Q vssd1 vssd1 vccd1 vccd1 hold3421/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4177 _17210_/Q vssd1 vssd1 vccd1 vccd1 hold4177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3432 _17241_/Q vssd1 vssd1 vccd1 vccd1 hold3432/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4188 _12142_/X vssd1 vssd1 vccd1 vccd1 _17204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3443 _12145_/X vssd1 vssd1 vccd1 vccd1 _17205_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3454 _17272_/Q vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4199 _15997_/Q vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2720 _08020_/X vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3465 _12037_/X vssd1 vssd1 vccd1 vccd1 _17169_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3476 _16745_/Q vssd1 vssd1 vccd1 vccd1 hold3476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2731 _15739_/Q vssd1 vssd1 vccd1 vccd1 hold2731/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2742 _08095_/X vssd1 vssd1 vccd1 vccd1 _15687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3487 _11482_/X vssd1 vssd1 vccd1 vccd1 _16984_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08988_ _15491_/A hold437/X vssd1 vssd1 vccd1 vccd1 _16111_/D sky130_fd_sc_hd__and2_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3498 _17367_/Q vssd1 vssd1 vccd1 vccd1 hold3498/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2753 _17957_/Q vssd1 vssd1 vccd1 vccd1 hold2753/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2764 _14103_/X vssd1 vssd1 vccd1 vccd1 _17854_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2775 _14673_/X vssd1 vssd1 vccd1 vccd1 _18127_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2786 _08016_/X vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07939_ _14735_/A hold203/X vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__or2_4
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2797 _16159_/Q vssd1 vssd1 vccd1 vccd1 hold2797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10950_ _11052_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _09987_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__or2_1
X_10881_ _11553_/A _10881_/B vssd1 vssd1 vccd1 vccd1 _10881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ hold3431/X _12619_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ hold3586/X _12550_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__mux2_1
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _12057_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12482_ _17334_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__or2_1
X_15270_ hold695/X _15486_/A2 _09357_/B hold536/X vssd1 vssd1 vccd1 vccd1 _15270_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14221_ hold1847/X _14216_/Y _14220_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14221_/X
+ sky130_fd_sc_hd__o211a_1
X_11433_ _12204_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14152_ _15551_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__or2_1
X_11364_ _12243_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ hold3972/X _10637_/B _10314_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10315_/X
+ sky130_fd_sc_hd__o211a_1
X_13103_ _13311_/A1 _13101_/X _13102_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14083_ hold1377/X _14094_/B _14082_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11295_ _12243_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13034_ hold960/X _13056_/C _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__and4_1
Xhold5390 _12127_/X vssd1 vssd1 vccd1 vccd1 _17199_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17911_ _18039_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
X_10246_ hold3718/X _10628_/B _10245_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10246_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17842_ _17842_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10177_ hold4897/X _10601_/B _10176_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17773_ _17871_/CLK _17773_/D vssd1 vssd1 vccd1 vccd1 _17773_/Q sky130_fd_sc_hd__dfxtp_1
X_14985_ hold3106/X _15004_/B _14984_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16724_ _18058_/CLK _16724_/D vssd1 vssd1 vccd1 vccd1 _16724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13936_ _14330_/A hold1291/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13937_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16655_ _18153_/CLK _16655_/D vssd1 vssd1 vccd1 vccd1 _16655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13867_ _13873_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _17742_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_187_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _17623_/CLK _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12818_ hold3187/X _12817_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12818_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_232_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16586_ _18142_/CLK _16586_/D vssd1 vssd1 vccd1 vccd1 _16586_/Q sky130_fd_sc_hd__dfxtp_1
X_13798_ hold3890/X _13798_/A2 _13797_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _13798_/X
+ sky130_fd_sc_hd__o211a_1
X_18325_ _18383_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _15537_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__or2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ hold3209/X _12748_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18256_ _18350_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15468_ hold667/X _09367_/A _15479_/B1 hold337/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17207_ _17207_/CLK _17207_/D vssd1 vssd1 vccd1 vccd1 _17207_/Q sky130_fd_sc_hd__dfxtp_1
X_14419_ _15099_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18187_ _18219_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15399_ hold714/X _09365_/B _09392_/C hold737/X _15398_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold604 hold604/A vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dlygate4sd3_1
X_17138_ _17170_/CLK _17138_/D vssd1 vssd1 vccd1 vccd1 _17138_/Q sky130_fd_sc_hd__dfxtp_1
Xhold615 hold615/A vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 hold626/A vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold637 hold637/A vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 hold648/A vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17069_ _17883_/CLK _17069_/D vssd1 vssd1 vccd1 vccd1 _17069_/Q sky130_fd_sc_hd__dfxtp_1
Xhold659 hold659/A vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08911_ _12424_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _16073_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09891_ _09963_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__or2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_398_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17898_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _08320_/X vssd1 vssd1 vccd1 vccd1 _15793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _07975_/X vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 _16219_/Q vssd1 vssd1 vccd1 vccd1 hold2027/X sky130_fd_sc_hd__dlygate4sd3_1
X_08842_ hold402/X hold672/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold673/A sky130_fd_sc_hd__mux2_1
Xhold2038 _15780_/Q vssd1 vssd1 vccd1 vccd1 hold2038/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1304 _08251_/X vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_327_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17871_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2049 _16153_/Q vssd1 vssd1 vccd1 vccd1 hold2049/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1315 _08061_/X vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 _09298_/X vssd1 vssd1 vccd1 vccd1 _16259_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1337 _14905_/X vssd1 vssd1 vccd1 vccd1 _18238_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ hold228/X hold422/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold423/A sky130_fd_sc_hd__mux2_1
Xhold1348 _17758_/Q vssd1 vssd1 vccd1 vccd1 hold1348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _17832_/Q vssd1 vssd1 vccd1 vccd1 hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ _15547_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _12738_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _16239_/D sky130_fd_sc_hd__and2_1
XFILLER_0_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ _14946_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17876_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09187_ hold2677/X _09218_/B _09186_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _09187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ hold246/A _15708_/Q hold240/X vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08069_ hold2357/X _08097_/A2 _08068_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10100_ hold1346/X hold4599/X _10580_/C vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ hold5515/X _11753_/B _11079_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3240 hold5855/X vssd1 vssd1 vccd1 vccd1 hold5856/A sky130_fd_sc_hd__buf_6
XTAP_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _10031_/A _10055_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__and3_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3251 _17487_/Q vssd1 vssd1 vccd1 vccd1 hold3251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3262 _16714_/Q vssd1 vssd1 vccd1 vccd1 hold3262/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3273 _17507_/Q vssd1 vssd1 vccd1 vccd1 hold3273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3284 _12959_/X vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3295 _16335_/Q vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2550 _17860_/Q vssd1 vssd1 vccd1 vccd1 hold2550/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2561 _07876_/X vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 _15701_/Q vssd1 vssd1 vccd1 vccd1 hold2572/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2583 _17958_/Q vssd1 vssd1 vccd1 vccd1 hold2583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2594 _17906_/Q vssd1 vssd1 vccd1 vccd1 hold2594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1860 _14779_/X vssd1 vssd1 vccd1 vccd1 _18178_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1871 hold6051/X vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__buf_1
X_14770_ _14878_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _12057_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__or2_1
Xhold1882 _09231_/X vssd1 vssd1 vccd1 vccd1 _16227_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1893 _18385_/Q vssd1 vssd1 vccd1 vccd1 hold1893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13721_ hold1793/X hold5709/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10933_ hold4539/X _11207_/B _10932_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _18319_/CLK _16440_/D vssd1 vssd1 vccd1 vccd1 _16440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ hold3806/X _11726_/B _10863_/X _12981_/A vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__o211a_1
X_13652_ hold1674/X _17671_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13653_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_49_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_49_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12603_ _13002_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _17377_/D sky130_fd_sc_hd__and2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _18346_/CLK _16371_/D vssd1 vssd1 vccd1 vccd1 _16371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ hold5042/X _11177_/B _10794_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10795_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ hold1192/X hold4297/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__mux2_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18110_ _18234_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15322_ _15489_/A _15322_/B _15322_/C _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/X
+ sky130_fd_sc_hd__or4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ _13002_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _17354_/D sky130_fd_sc_hd__and2_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18041_ _18041_/CLK hold798/X vssd1 vssd1 vccd1 vccd1 hold797/A sky130_fd_sc_hd__dfxtp_1
X_15253_ _15490_/A1 _15245_/X _15252_/X _15490_/B1 hold5854/A vssd1 vssd1 vccd1 vccd1
+ _15253_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ hold65/X _12509_/A2 _12507_/A3 _12464_/X _15364_/A vssd1 vssd1 vccd1 vccd1
+ hold66/A sky130_fd_sc_hd__o311a_1
XFILLER_0_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14204_ _14328_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ hold4495/X _12344_/B _11415_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11416_/X
+ sky130_fd_sc_hd__o211a_1
X_15184_ hold1811/X _15219_/B _15183_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15184_/X
+ sky130_fd_sc_hd__o211a_1
X_12396_ _12396_/A hold779/X vssd1 vssd1 vccd1 vccd1 _17291_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ hold1527/X _14142_/B _14134_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _14135_/X
+ sky130_fd_sc_hd__o211a_1
X_11347_ hold4103/X _11729_/B _11346_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_238_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14066_ _14854_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14066_/X sky130_fd_sc_hd__or2_1
X_11278_ hold5555/X _11762_/B _11277_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11278_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10229_ hold1954/X hold3752/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__mux2_1
X_13017_ _14910_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_420_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17253_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17825_ _17825_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _17852_/CLK _17756_/D vssd1 vssd1 vccd1 vccd1 _17756_/Q sky130_fd_sc_hd__dfxtp_1
X_14968_ _14968_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16707_ _18216_/CLK _16707_/D vssd1 vssd1 vccd1 vccd1 _16707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13919_ _13919_/A _13919_/B vssd1 vssd1 vccd1 vccd1 _17765_/D sky130_fd_sc_hd__and2_1
XFILLER_0_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17687_ _17693_/CLK _17687_/D vssd1 vssd1 vccd1 vccd1 _17687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14899_ hold1875/X _14896_/Y _14898_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638_ _18182_/CLK _16638_/D vssd1 vssd1 vccd1 vccd1 _16638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16569_ _18163_/CLK _16569_/D vssd1 vssd1 vccd1 vccd1 _16569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ _15551_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__or2_1
X_18308_ _18396_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09041_ _12438_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _16137_/D sky130_fd_sc_hd__and2_1
X_18239_ _18413_/CLK hold941/X vssd1 vssd1 vccd1 vccd1 hold940/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold401 input15/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__buf_1
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold412 hold412/A vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 hold423/A vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold434 hold434/A vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold445 hold466/X vssd1 vssd1 vccd1 vccd1 hold467/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold456 hold456/A vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold467 hold467/A vssd1 vssd1 vccd1 vccd1 input44/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold489 hold489/A vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ hold4831/X _10055_/B _09942_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09943_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout903 _14894_/A vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__buf_8
XFILLER_0_106_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout914 _15173_/A vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout925 hold998/X vssd1 vssd1 vccd1 vccd1 hold915/A sky130_fd_sc_hd__buf_6
XFILLER_0_42_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout936 _15207_/A vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09874_ hold5226/X _10070_/B _09873_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_161_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18303_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout947 hold1152/X vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__buf_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _15520_/X vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 hold1112/A vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08825_ _15364_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _16031_/D sky130_fd_sc_hd__and2_1
Xhold1123 _16156_/Q vssd1 vssd1 vccd1 vccd1 hold1123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 la_data_in[15] vssd1 vssd1 vccd1 vccd1 hold1134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 _15849_/Q vssd1 vssd1 vccd1 vccd1 hold1145/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 input52/X vssd1 vssd1 vccd1 vccd1 hold1156/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1167 _09195_/X vssd1 vssd1 vccd1 vccd1 _16209_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _15414_/A hold272/X vssd1 vssd1 vccd1 vccd1 _15998_/D sky130_fd_sc_hd__and2_1
Xhold1178 _18315_/Q vssd1 vssd1 vccd1 vccd1 hold1178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _08516_/X vssd1 vssd1 vccd1 vccd1 _15885_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ hold361/X hold649/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold650/A sky130_fd_sc_hd__mux2_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09308_ hold3002/X _09325_/B _09307_/X _12600_/A vssd1 vssd1 vccd1 vccd1 _09308_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ _16684_/Q _10598_/B _10580_/C vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09239_ _15515_/A hold2765/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _12344_/A _12274_/A2 _12249_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11201_ _16891_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__and3_1
XFILLER_0_146_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ hold4451/X _13877_/B _12180_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_249_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18198_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11132_ hold2943/X _16868_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _11133_/B sky130_fd_sc_hd__mux2_1
Xhold990 hold990/A vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__clkbuf_4
X_15940_ _17314_/CLK _15940_/D vssd1 vssd1 vccd1 vccd1 hold617/A sky130_fd_sc_hd__dfxtp_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ hold1781/X hold5066/X _11159_/C vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3070 _14424_/X vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10014_ _13150_/A _09918_/A _10013_/X vssd1 vssd1 vccd1 vccd1 _10014_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3081 _14416_/X vssd1 vssd1 vccd1 vccd1 _18004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3092 _18302_/Q vssd1 vssd1 vccd1 vccd1 hold3092/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _17742_/CLK _15871_/D vssd1 vssd1 vccd1 vccd1 _15871_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 _18135_/Q vssd1 vssd1 vccd1 vccd1 hold2380/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _17745_/CLK _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14822_ _15215_/A _14826_/B vssd1 vssd1 vccd1 vccd1 _14822_/Y sky130_fd_sc_hd__nand2_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2391 _15766_/Q vssd1 vssd1 vccd1 vccd1 hold2391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _18384_/CLK _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _15098_/X vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14753_ hold3122/X _14774_/B _14752_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14753_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11965_ hold4263/X _12347_/B _11964_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13800_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ hold3118/X _16796_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17472_ _17879_/CLK _17472_/D vssd1 vssd1 vccd1 vccd1 _17472_/Q sky130_fd_sc_hd__dfxtp_1
X_14684_ _15131_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ hold4085/X _12374_/B _11895_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11896_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16423_ _18366_/CLK _16423_/D vssd1 vssd1 vccd1 vccd1 _16423_/Q sky130_fd_sc_hd__dfxtp_1
X_13635_ _13767_/A _13635_/B vssd1 vssd1 vccd1 vccd1 _13635_/X sky130_fd_sc_hd__or2_1
X_10847_ hold2818/X hold5481/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16354_ _18265_/CLK _16354_/D vssd1 vssd1 vccd1 vccd1 _16354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _13788_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__or2_1
X_10778_ hold3222/X _16750_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15305_ hold814/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12517_ hold1179/X hold3153/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16285_ _18459_/CLK _16285_/D vssd1 vssd1 vccd1 vccd1 _16285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13791_/A _13497_/B vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__or2_1
X_18024_ _18124_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
X_15236_ _17327_/Q _15448_/B1 _15485_/B1 hold480/X vssd1 vssd1 vccd1 vccd1 _15236_/X
+ sky130_fd_sc_hd__a22o_1
X_12448_ _17317_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15167_ _15547_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15167_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12379_ _13888_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _17283_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_240_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14118_ _14403_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ hold1689/X _15113_/B _15097_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15098_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14049_ hold2276/X _14038_/B _14048_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _09061_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _15927_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09590_ hold1857/X _13302_/A _10580_/C vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__mux2_1
X_17808_ _17808_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08541_ _12438_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _15894_/D sky130_fd_sc_hd__and2_1
X_17739_ _17739_/CLK _17739_/D vssd1 vssd1 vccd1 vccd1 _17739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08472_ _14758_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ hold271/X hold647/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__mux2_1
Xhold5901 _13056_/C vssd1 vssd1 vccd1 vccd1 hold5901/X sky130_fd_sc_hd__buf_1
XFILLER_0_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5912 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold5912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5923 _17537_/Q vssd1 vssd1 vccd1 vccd1 hold5923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5934 _17539_/Q vssd1 vssd1 vccd1 vccd1 hold5934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 hold13/X vssd1 vssd1 vccd1 vccd1 input22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5945 _17530_/Q vssd1 vssd1 vccd1 vccd1 hold5945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5956 data_in[12] vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_342_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17585_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5967 data_in[30] vssd1 vssd1 vccd1 vccd1 hold495/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5978 _17947_/Q vssd1 vssd1 vccd1 vccd1 hold5978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5989 _18352_/Q vssd1 vssd1 vccd1 vccd1 hold5989/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _12396_/A vssd1 vssd1 vccd1 vccd1 _12386_/A sky130_fd_sc_hd__clkbuf_4
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout711 _13037_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09926_ hold3008/X _16466_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__mux2_1
Xfanout722 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _14434_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout733 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout744 _08377_/A vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__buf_4
Xfanout755 _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__buf_4
Xfanout766 _14538_/C1 vssd1 vssd1 vccd1 vccd1 _14131_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09857_ hold1996/X _16443_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout777 _08349_/A vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__buf_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 fanout796/X vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_225_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout799 _09976_/C1 vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ hold215/X hold337/X _08808_/S vssd1 vssd1 vccd1 vccd1 hold338/A sky130_fd_sc_hd__mux2_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ hold1689/X _16420_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ hold88/X hold90/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__mux2_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _17074_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ _11100_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__or2_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ hold2735/X hold4982/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13420_ hold4171/X _13802_/B _13419_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13420_/X
+ sky130_fd_sc_hd__o211a_1
X_10632_ hold4639/X _10536_/A _10631_/X vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__or2_1
X_13351_ hold5695/X _13829_/B _13350_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _17258_/Q _13811_/B _12302_/C vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__and3_1
X_16070_ _16077_/CLK _16070_/D vssd1 vssd1 vccd1 vccd1 _16070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10554_/A _10494_/B vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__or2_1
X_13282_ _17586_/Q _17120_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ _15183_/A hold1601/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15021_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ hold2248/X hold5308/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__mux2_1
X_12164_ hold2343/X hold5364/X _13862_/C vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__mux2_1
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12095_ hold2743/X hold3918/X _13412_/S vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__mux2_1
X_16972_ _17882_/CLK _16972_/D vssd1 vssd1 vccd1 vccd1 _16972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15923_ _16087_/CLK _15923_/D vssd1 vssd1 vccd1 vccd1 hold893/A sky130_fd_sc_hd__dfxtp_1
X_11046_ _11052_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/X sky130_fd_sc_hd__or2_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _17613_/CLK _15854_/D vssd1 vssd1 vccd1 vccd1 _15854_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ hold1829/X _14828_/B _14804_/X _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14805_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _17748_/CLK _15785_/D vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ hold1385/X _17510_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17524_ _17525_/CLK hold934/X vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_176_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _15183_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__or2_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11948_ hold2428/X hold4087/X _13868_/C vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17455_ _17455_/CLK _17455_/D vssd1 vssd1 vccd1 vccd1 _17455_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ hold2687/X _14666_/B _14666_/Y _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14667_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11879_ _15709_/Q hold3625/X _12362_/C vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__mux2_1
X_16406_ _18349_/CLK _16406_/D vssd1 vssd1 vccd1 vccd1 _16406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ hold3428/X _13808_/B _13617_/X _12657_/A vssd1 vssd1 vccd1 vccd1 _13618_/X
+ sky130_fd_sc_hd__o211a_1
X_17386_ _18435_/CLK _17386_/D vssd1 vssd1 vccd1 vccd1 _17386_/Q sky130_fd_sc_hd__dfxtp_1
X_14598_ _15099_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ _18376_/CLK _16337_/D vssd1 vssd1 vccd1 vccd1 _16337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ hold4559/X _13856_/B _13548_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16268_ _17370_/CLK _16268_/D vssd1 vssd1 vccd1 vccd1 _16268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5208 _16945_/Q vssd1 vssd1 vccd1 vccd1 hold5208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5219 _12022_/X vssd1 vssd1 vccd1 vccd1 _17164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _18429_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_207_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4507 _17744_/Q vssd1 vssd1 vccd1 vccd1 hold4507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4518 _12085_/X vssd1 vssd1 vccd1 vccd1 _17185_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16199_ _17479_/CLK _16199_/D vssd1 vssd1 vccd1 vccd1 _16199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4529 _17271_/Q vssd1 vssd1 vccd1 vccd1 hold4529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3806 _16810_/Q vssd1 vssd1 vccd1 vccd1 hold3806/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3817 _16623_/Q vssd1 vssd1 vccd1 vccd1 hold3817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3828 _09835_/X vssd1 vssd1 vccd1 vccd1 _16435_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3839 _16568_/Q vssd1 vssd1 vccd1 vccd1 hold3839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07972_ _15541_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ _11064_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09984_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09573_ _10467_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08524_ hold554/X hold790/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold791/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08455_ hold2672/X _08488_/B _08454_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08386_ _14782_/A hold2194/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ _09061_/A hold282/X vssd1 vssd1 vccd1 vccd1 _16120_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5720 _13576_/X vssd1 vssd1 vccd1 vccd1 _17645_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5731 _17667_/Q vssd1 vssd1 vccd1 vccd1 hold5731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5742 _13540_/X vssd1 vssd1 vccd1 vccd1 _17633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5753 _17601_/Q vssd1 vssd1 vccd1 vccd1 hold5753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5764 output88/X vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_12
Xhold5775 hold5928/X vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5786 hold5786/A vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_12
Xhold5797 hold5937/X vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout530 _09166_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__buf_4
Xfanout541 _08486_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__buf_6
X_09909_ _09987_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__or2_1
Xfanout552 _08268_/B vssd1 vssd1 vccd1 vccd1 _08263_/A2 sky130_fd_sc_hd__buf_8
Xfanout563 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08029_/B sky130_fd_sc_hd__buf_8
Xfanout574 _14602_/B vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout585 _13305_/B vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__buf_4
XFILLER_0_191_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ hold3322/X _12919_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__mux2_1
Xfanout596 _12985_/S vssd1 vssd1 vccd1 vccd1 _12922_/S sky130_fd_sc_hd__buf_6
XFILLER_0_226_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ hold3421/X _12850_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11802_ hold3862/X _12246_/A _11801_/X vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _17145_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ hold3342/X _12781_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14521_ _15201_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14521_/X sky130_fd_sc_hd__or2_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ hold4751/X _11553_/A _11732_/X vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__a21oi_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17269_/CLK _17240_/D vssd1 vssd1 vccd1 vccd1 _17240_/Q sky130_fd_sc_hd__dfxtp_1
X_14452_ hold1263/X _14482_/A2 _14451_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14452_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ _11670_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ hold2439/X hold3641/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10615_ _18461_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _16695_/D sky130_fd_sc_hd__nor2_1
X_17171_ _17171_/CLK _17171_/D vssd1 vssd1 vccd1 vccd1 _17171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_264_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18059_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14383_ _14330_/A hold1129/X hold333/X vssd1 vssd1 vccd1 vccd1 _14384_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11595_ _12243_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16122_ _16127_/CLK _16122_/D vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13334_ hold1312/X _17565_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__mux2_1
X_10546_ hold4008/X _10646_/B _10545_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16053_ _16089_/CLK _16053_/D vssd1 vssd1 vccd1 vccd1 hold661/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13265_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__and2_1
X_10477_ _10571_/A _10477_/A2 _10476_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10477_/X
+ sky130_fd_sc_hd__o211a_1
X_15004_ _15004_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_161_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12216_ _12261_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__or2_1
X_13196_ hold4678/X _13195_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12147_ _12243_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12078_ _13461_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__or2_1
X_16955_ _17821_/CLK _16955_/D vssd1 vssd1 vccd1 vccd1 _16955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15906_ _17315_/CLK _15906_/D vssd1 vssd1 vccd1 vccd1 hold519/A sky130_fd_sc_hd__dfxtp_1
X_11029_ hold4531/X _11207_/B _11028_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11029_/X
+ sky130_fd_sc_hd__o211a_1
X_16886_ _18026_/CLK _16886_/D vssd1 vssd1 vccd1 vccd1 _16886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_8_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_15837_ _17696_/CLK _15837_/D vssd1 vssd1 vccd1 vccd1 _15837_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ _17693_/CLK _15768_/D vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14719_ hold1941/X _14714_/B _14718_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14719_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17507_ _17507_/CLK _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15699_ _17899_/CLK _15699_/D vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08240_ _14854_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08240_/X sky130_fd_sc_hd__or2_1
X_17438_ _18434_/CLK _17438_/D vssd1 vssd1 vccd1 vccd1 _17438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_15 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _08759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_37 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _12804_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _15723_/D sky130_fd_sc_hd__and2_1
X_17369_ _17370_/CLK _17369_/D vssd1 vssd1 vccd1 vccd1 _17369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_59 hold746/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5005 _11769_/Y vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5016 _16755_/Q vssd1 vssd1 vccd1 vccd1 hold5016/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5027 _10444_/X vssd1 vssd1 vccd1 vccd1 _16638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput100 _13105_/A vssd1 vssd1 vccd1 vccd1 hold5786/A sky130_fd_sc_hd__buf_6
Xhold5038 _16440_/Q vssd1 vssd1 vccd1 vccd1 hold5038/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5049 _09700_/X vssd1 vssd1 vccd1 vccd1 _16390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput111 hold5890/X vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_12
Xhold4304 _13495_/X vssd1 vssd1 vccd1 vccd1 _17618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4315 _17673_/Q vssd1 vssd1 vccd1 vccd1 hold4315/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput122 hold5888/X vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput133 hold5837/X vssd1 vssd1 vccd1 vccd1 hold5838/A sky130_fd_sc_hd__buf_6
Xhold4326 _11317_/X vssd1 vssd1 vccd1 vccd1 _16929_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4337 _10759_/X vssd1 vssd1 vccd1 vccd1 _16743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput144 hold5862/X vssd1 vssd1 vccd1 vccd1 load_status[4] sky130_fd_sc_hd__buf_12
Xhold3603 _12351_/Y vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4348 _17638_/Q vssd1 vssd1 vccd1 vccd1 hold4348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3614 _09679_/X vssd1 vssd1 vccd1 vccd1 _16383_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4359 _13552_/X vssd1 vssd1 vccd1 vccd1 _17637_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3625 _17117_/Q vssd1 vssd1 vccd1 vccd1 hold3625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3636 _09667_/X vssd1 vssd1 vccd1 vccd1 _16379_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2902 _09294_/X vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3647 _17579_/Q vssd1 vssd1 vccd1 vccd1 hold3647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2913 _18454_/Q vssd1 vssd1 vccd1 vccd1 hold2913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3658 _09781_/X vssd1 vssd1 vccd1 vccd1 _16417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3669 _10312_/X vssd1 vssd1 vccd1 vccd1 _16594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 _09155_/X vssd1 vssd1 vccd1 vccd1 _16190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2935 _18195_/Q vssd1 vssd1 vccd1 vccd1 hold2935/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18405_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2946 _08196_/X vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07955_ hold1684/X _07991_/A2 _07954_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07955_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2957 _17948_/Q vssd1 vssd1 vccd1 vccd1 hold2957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 _14865_/X vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2979 _18334_/Q vssd1 vssd1 vccd1 vccd1 hold2979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07886_ _15509_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ hold3405/X _10025_/B _09624_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09625_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09556_ hold4759/X _10034_/B _09555_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ hold999/X _08517_/B vssd1 vssd1 vccd1 vccd1 _08507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09487_ _13056_/C _13029_/A _13034_/D hold960/X vssd1 vssd1 vccd1 vccd1 _13035_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08438_ hold1145/X _08440_/A2 _08437_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ _08369_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _15816_/D sky130_fd_sc_hd__and2_1
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10400_ hold2353/X _16624_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ hold5453/X _11762_/B _11379_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11380_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ hold1952/X _16601_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5550 _10732_/X vssd1 vssd1 vccd1 vccd1 _16734_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13050_ hold5859/X hold960/X _13055_/C vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__a21o_2
X_10262_ hold3075/X hold4042/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10263_/B sky130_fd_sc_hd__mux2_1
Xhold5561 _16981_/Q vssd1 vssd1 vccd1 vccd1 hold5561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5572 _09544_/X vssd1 vssd1 vccd1 vccd1 _16338_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5583 _16869_/Q vssd1 vssd1 vccd1 vccd1 hold5583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5594 _11107_/X vssd1 vssd1 vccd1 vccd1 _16859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12001_ hold3918/X _12293_/B _12000_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4860 _10288_/X vssd1 vssd1 vccd1 vccd1 _16586_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10193_ hold2750/X hold3689/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__mux2_1
Xhold4871 _17105_/Q vssd1 vssd1 vccd1 vccd1 hold4871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4882 _11196_/Y vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4893 _16889_/Q vssd1 vssd1 vccd1 vccd1 hold4893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout360 _15211_/B vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__buf_6
Xfanout371 _15016_/B vssd1 vssd1 vccd1 vccd1 _15018_/B sky130_fd_sc_hd__buf_6
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout382 _14788_/Y vssd1 vssd1 vccd1 vccd1 _14826_/B sky130_fd_sc_hd__buf_6
X_16740_ _18049_/CLK _16740_/D vssd1 vssd1 vccd1 vccd1 _16740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13952_ _15513_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13952_/X sky130_fd_sc_hd__or2_1
Xfanout393 _14535_/B vssd1 vssd1 vccd1 vccd1 _14541_/B sky130_fd_sc_hd__buf_6
XFILLER_0_205_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ _12909_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _17477_/D sky130_fd_sc_hd__and2_1
X_16671_ _18227_/CLK _16671_/D vssd1 vssd1 vccd1 vccd1 _16671_/Q sky130_fd_sc_hd__dfxtp_1
X_13883_ _17748_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__and3_1
XFILLER_0_213_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18410_ _18410_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15622_ _17274_/CLK _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _12912_/A _12834_/B vssd1 vssd1 vccd1 vccd1 _17454_/D sky130_fd_sc_hd__and2_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18341_/CLK hold561/X vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12765_ _12768_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _17431_/D sky130_fd_sc_hd__and2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_445_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17254_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14504_ hold1781/X _14535_/B _14503_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14504_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _18272_/CLK hold939/X vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ hold5106/X _12308_/B _11715_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11716_/X
+ sky130_fd_sc_hd__o211a_1
X_15484_ hold363/X _15484_/A2 _15484_/B1 hold519/X vssd1 vssd1 vccd1 vccd1 _15489_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _17408_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ _17444_/CLK _17223_/D vssd1 vssd1 vccd1 vccd1 _17223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14435_ _15169_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11647_ hold5242/X _11747_/B _11646_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11647_/X
+ sky130_fd_sc_hd__o211a_1
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_6
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 input24/A vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_6
X_17154_ _17237_/CLK _17154_/D vssd1 vssd1 vccd1 vccd1 _17154_/Q sky130_fd_sc_hd__dfxtp_1
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
X_14366_ _14366_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _17980_/D sky130_fd_sc_hd__and2_1
Xinput46 input46/A vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
X_11578_ hold4360/X _11584_/A2 _11577_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11578_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
X_16105_ _17340_/CLK _16105_/D vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput68 input68/A vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_13317_ _13797_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold808 hold808/A vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__buf_6
Xhold819 hold824/X vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__clkbuf_4
X_10529_ hold1887/X hold4811/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10530_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17085_ _17863_/CLK _17085_/D vssd1 vssd1 vccd1 vccd1 _17085_/Q sky130_fd_sc_hd__dfxtp_1
X_14297_ hold1003/X hold756/X _14296_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _14297_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _17327_/CLK _16036_/D vssd1 vssd1 vccd1 vccd1 hold434/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _13241_/X _13247_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _13178_/X hold5919/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__mux2_1
Xhold2209 _15084_/X vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1508 _13908_/X vssd1 vssd1 vccd1 vccd1 _13909_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ _18019_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 hold658/A sky130_fd_sc_hd__dfxtp_1
Xhold1519 _18230_/Q vssd1 vssd1 vccd1 vccd1 hold1519/X sky130_fd_sc_hd__dlygate4sd3_1
X_16938_ _17816_/CLK _16938_/D vssd1 vssd1 vccd1 vccd1 _16938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16869_ _18070_/CLK _16869_/D vssd1 vssd1 vccd1 vccd1 _16869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09410_ _09438_/B _16291_/Q vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09341_ _18458_/Q _07802_/B _15490_/A1 vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_133_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_186_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09272_ _12747_/A hold535/X vssd1 vssd1 vccd1 vccd1 _16247_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17329_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08223_ _15557_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _15559_/A hold1737/X hold240/X vssd1 vssd1 vccd1 vccd1 _08154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08085_ hold2107/X _08088_/B _08084_/Y _08127_/A vssd1 vssd1 vccd1 vccd1 _08085_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4101 _17624_/Q vssd1 vssd1 vccd1 vccd1 hold4101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4112 _16015_/Q vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4123 _16388_/Q vssd1 vssd1 vccd1 vccd1 hold4123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4134 _13321_/X vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3400 _09613_/X vssd1 vssd1 vccd1 vccd1 _16361_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4145 _17171_/Q vssd1 vssd1 vccd1 vccd1 hold4145/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4156 _11134_/X vssd1 vssd1 vccd1 vccd1 _16868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3411 _12716_/X vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3422 _16363_/Q vssd1 vssd1 vccd1 vccd1 hold3422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4167 _13519_/X vssd1 vssd1 vccd1 vccd1 _17626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4178 _12064_/X vssd1 vssd1 vccd1 vccd1 _17178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3433 _12157_/X vssd1 vssd1 vccd1 vccd1 _17209_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3444 _16838_/Q vssd1 vssd1 vccd1 vccd1 hold3444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4189 _16868_/Q vssd1 vssd1 vccd1 vccd1 hold4189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2710 _14333_/X vssd1 vssd1 vccd1 vccd1 _17964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3455 _12250_/X vssd1 vssd1 vccd1 vccd1 _17240_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2721 _18025_/Q vssd1 vssd1 vccd1 vccd1 hold2721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3466 _17396_/Q vssd1 vssd1 vccd1 vccd1 hold3466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2732 _08206_/X vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08987_ hold210/X hold436/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold437/A sky130_fd_sc_hd__mux2_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3477 _10669_/X vssd1 vssd1 vccd1 vccd1 _16713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3488 _17366_/Q vssd1 vssd1 vccd1 vccd1 hold3488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _15625_/Q vssd1 vssd1 vccd1 vccd1 hold2743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3499 _12572_/X vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2754 _14319_/X vssd1 vssd1 vccd1 vccd1 _17957_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2765 _16231_/Q vssd1 vssd1 vccd1 vccd1 hold2765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _14735_/A hold203/X vssd1 vssd1 vccd1 vccd1 _07938_/Y sky130_fd_sc_hd__nor2_1
Xhold2776 _17853_/Q vssd1 vssd1 vccd1 vccd1 hold2776/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2787 _18130_/Q vssd1 vssd1 vccd1 vccd1 hold2787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2798 _09089_/X vssd1 vssd1 vccd1 vccd1 _16159_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07869_ _14774_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09608_ hold1479/X hold3860/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _17985_/Q hold4215/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10881_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_39_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_39_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ hold1070/X _13166_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__mux2_1
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ hold1325/X _17361_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ hold2293/X hold3523/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__mux2_1
X_12481_ hold53/X _12445_/A _12445_/B _12480_/X _12436_/A vssd1 vssd1 vccd1 vccd1
+ hold54/A sky130_fd_sc_hd__o311a_1
XFILLER_0_124_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14220_ _15185_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14220_/X sky130_fd_sc_hd__or2_1
X_11432_ hold993/X hold3932/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ hold2312/X _14148_/B _14150_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _14151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11363_ hold1712/X _16945_/Q _11594_/S vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ _13102_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _10542_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14082_ _15535_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14082_/X sky130_fd_sc_hd__or2_1
X_11294_ _17768_/Q hold3722/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5380 _10723_/X vssd1 vssd1 vccd1 vccd1 _16731_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13033_ _13056_/C hold922/X _13032_/Y vssd1 vssd1 vccd1 vccd1 hold923/A sky130_fd_sc_hd__a21oi_1
X_17910_ _18070_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _10497_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__or2_1
Xhold5391 _17134_/Q vssd1 vssd1 vccd1 vccd1 hold5391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4690 _11778_/Y vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _10488_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
X_17841_ _17871_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14984_ _14984_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__or2_1
X_17772_ _17899_/CLK hold276/X vssd1 vssd1 vccd1 vccd1 _17772_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout190 _13886_/B vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__buf_4
X_16723_ _18319_/CLK _16723_/D vssd1 vssd1 vccd1 vccd1 _16723_/Q sky130_fd_sc_hd__dfxtp_1
X_13935_ _13935_/A _13935_/B vssd1 vssd1 vccd1 vccd1 _17773_/D sky130_fd_sc_hd__and2_1
XFILLER_0_96_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ _18210_/CLK _16654_/D vssd1 vssd1 vccd1 vccd1 _16654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13866_ hold4012/X _12267_/A _13865_/X vssd1 vssd1 vccd1 vccd1 _13866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15605_ _17221_/CLK _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
X_12817_ hold2401/X _17450_/Q _12826_/S vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__mux2_1
X_16585_ _18141_/CLK _16585_/D vssd1 vssd1 vccd1 vccd1 _16585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13797_ _13797_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18324_ _18350_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_15536_ hold1499/X _15547_/B _15535_/X _12657_/A vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _16247_/Q _17427_/Q _12748_/S vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18255_ _18293_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ hold440/X _09365_/B _09362_/D _16127_/Q vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12679_ hold2632/X hold3756/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17206_ _17270_/CLK _17206_/D vssd1 vssd1 vccd1 vccd1 _17206_/Q sky130_fd_sc_hd__dfxtp_1
X_14418_ hold1267/X _14433_/B _14417_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _14418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18186_ _18186_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ hold699/X _09386_/A _15451_/A2 hold780/X vssd1 vssd1 vccd1 vccd1 _15398_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _17265_/CLK _17137_/D vssd1 vssd1 vccd1 vccd1 _17137_/Q sky130_fd_sc_hd__dfxtp_1
X_14349_ _14403_/A hold2112/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold605 hold31/X vssd1 vssd1 vccd1 vccd1 input19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 hold616/A vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 hold627/A vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold649 hold649/A vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ _17822_/CLK _17068_/D vssd1 vssd1 vccd1 vccd1 _17068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _17315_/CLK _16019_/D vssd1 vssd1 vccd1 vccd1 hold584/A sky130_fd_sc_hd__dfxtp_1
X_08910_ hold353/X hold758/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09890_ hold2416/X hold5040/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2006 _18076_/Q vssd1 vssd1 vccd1 vccd1 hold2006/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08841_ _12404_/A _08841_/B vssd1 vssd1 vccd1 vccd1 _16039_/D sky130_fd_sc_hd__and2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _15656_/Q vssd1 vssd1 vccd1 vccd1 hold2017/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _09215_/X vssd1 vssd1 vccd1 vccd1 _16219_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2039 _08294_/X vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _15725_/Q vssd1 vssd1 vccd1 vccd1 hold1305/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _15698_/Q vssd1 vssd1 vccd1 vccd1 hold1316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 _16255_/Q vssd1 vssd1 vccd1 vccd1 hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ _15374_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _16006_/D sky130_fd_sc_hd__and2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1338 _18158_/Q vssd1 vssd1 vccd1 vccd1 hold1338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1349 _17766_/Q vssd1 vssd1 vccd1 vccd1 hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_367_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17736_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09324_ hold905/X _09325_/B _09323_/Y _12969_/A vssd1 vssd1 vccd1 vccd1 hold906/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09255_ _15531_/A hold2205/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08206_ hold2731/X _08209_/B _08205_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08206_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09186_ _15515_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08137_ _08137_/A hold591/X vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__and2_1
XFILLER_0_222_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17510_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_226_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _14862_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3230 _17374_/Q vssd1 vssd1 vccd1 vccd1 hold3230/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _10603_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _16500_/D sky130_fd_sc_hd__nor2_1
Xhold3241 _09391_/X vssd1 vssd1 vccd1 vccd1 _16283_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3252 _12932_/X vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3263 _11151_/Y vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3274 _17355_/Q vssd1 vssd1 vccd1 vccd1 hold3274/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3285 _17348_/Q vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__buf_2
Xhold2540 _17875_/Q vssd1 vssd1 vccd1 vccd1 hold2540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3296 _10014_/Y vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2551 _14117_/X vssd1 vssd1 vccd1 vccd1 _17860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2562 _16204_/Q vssd1 vssd1 vccd1 vccd1 hold2562/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 _17827_/Q vssd1 vssd1 vccd1 vccd1 hold2573/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2584 _14321_/X vssd1 vssd1 vccd1 vccd1 _17958_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1850 _09429_/X vssd1 vssd1 vccd1 vccd1 _16300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 _14211_/X vssd1 vssd1 vccd1 vccd1 _17906_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1861 _17881_/Q vssd1 vssd1 vccd1 vccd1 hold1861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1872 _09427_/X vssd1 vssd1 vccd1 vccd1 _16299_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11981_ hold1767/X _17151_/Q _12344_/C vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__mux2_1
Xhold1883 _17944_/Q vssd1 vssd1 vccd1 vccd1 hold1883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1894 _15210_/X vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ _13814_/A _13814_/B _13719_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _17693_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _11670_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10932_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ hold4352/X _13847_/B _13650_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13651_/X
+ sky130_fd_sc_hd__o211a_1
X_10863_ _11631_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ hold3286/X _12601_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _18351_/CLK _16370_/D vssd1 vssd1 vccd1 vccd1 _16370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13582_ hold4499/X _13847_/B _13581_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _13582_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _11082_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__or2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15321_ _16296_/Q _15477_/A2 _15487_/B1 hold580/X _15320_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/D sky130_fd_sc_hd__a221o_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12533_ hold3281/X _12532_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__mux2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18040_ _18040_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _15489_/A _15252_/B _15252_/C _15252_/D vssd1 vssd1 vccd1 vccd1 _15252_/X
+ sky130_fd_sc_hd__or4_1
X_12464_ _17325_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14203_ hold2624/X _14202_/B _14202_/Y _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14203_/X
+ sky130_fd_sc_hd__o211a_1
X_11415_ _12057_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__or2_1
X_15183_ _15183_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12395_ hold596/X hold778/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold779/A sky130_fd_sc_hd__mux2_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _15207_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14134_/X sky130_fd_sc_hd__or2_1
X_11346_ _11637_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__or2_1
XFILLER_0_240_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ hold2236/X _14107_/A2 _14064_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _14065_/X
+ sky130_fd_sc_hd__o211a_1
X_11277_ _11667_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11277_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13016_ hold1197/X _13003_/Y _13015_/X _12531_/A vssd1 vssd1 vccd1 vccd1 _13016_/X
+ sky130_fd_sc_hd__o211a_1
X_10228_ hold3744/X _10628_/B _10227_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _17884_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__buf_4
XFILLER_0_234_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ hold3728/X _10631_/B _10158_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_234_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14967_ hold754/X hold393/X vssd1 vssd1 vccd1 vccd1 _15016_/B sky130_fd_sc_hd__or2_4
X_17755_ _17883_/CLK _17755_/D vssd1 vssd1 vccd1 vccd1 _17755_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_460_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18442_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_222_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ _18198_/CLK _16706_/D vssd1 vssd1 vccd1 vccd1 _16706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13918_ _15207_/A hold1429/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__mux2_1
X_14898_ _14968_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__or2_1
X_17686_ _17686_/CLK _17686_/D vssd1 vssd1 vccd1 vccd1 _17686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16637_ _18225_/CLK _16637_/D vssd1 vssd1 vccd1 vccd1 _16637_/Q sky130_fd_sc_hd__dfxtp_1
X_13849_ _13873_/A _13849_/B vssd1 vssd1 vccd1 vccd1 _17736_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_202_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16568_ _17968_/CLK _16568_/D vssd1 vssd1 vccd1 vccd1 _16568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ _18309_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15519_ _15519_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__or2_1
X_16499_ _18384_/CLK _16499_/D vssd1 vssd1 vccd1 vccd1 _16499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09040_ hold353/X hold428/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18238_ _18367_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ _18201_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold402 hold44/X vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__buf_4
XFILLER_0_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold413 hold413/A vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold446 hold468/X vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__buf_6
XFILLER_0_29_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 input44/X vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _09960_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__or2_1
Xhold479 hold479/A vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout904 hold808/X vssd1 vssd1 vccd1 vccd1 _14894_/A sky130_fd_sc_hd__buf_8
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout915 hold1066/X vssd1 vssd1 vccd1 vccd1 hold1067/A sky130_fd_sc_hd__buf_4
Xfanout926 hold998/X vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__buf_4
X_09873_ _10191_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__or2_1
Xfanout937 _15207_/A vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__buf_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 hold1152/X vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__clkbuf_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ hold98/X hold768/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__mux2_1
Xhold1102 _18339_/Q vssd1 vssd1 vccd1 vccd1 hold1102/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1113 _09068_/X vssd1 vssd1 vccd1 vccd1 hold1113/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1124 _09083_/X vssd1 vssd1 vccd1 vccd1 _16156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 hold1135/A vssd1 vssd1 vccd1 vccd1 input43/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1146 _08438_/X vssd1 vssd1 vccd1 vccd1 _15849_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ hold271/X _15998_/Q _08779_/S vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__mux2_1
Xhold1157 _09400_/B vssd1 vssd1 vccd1 vccd1 _09122_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _18284_/Q vssd1 vssd1 vccd1 vccd1 hold1168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _17512_/Q vssd1 vssd1 vccd1 vccd1 hold1179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _09055_/A hold782/X vssd1 vssd1 vccd1 vccd1 _15964_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_130_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_240_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ _14988_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ _12768_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _16230_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ hold1521/X _09177_/A2 _09168_/X _12909_/A vssd1 vssd1 vccd1 vccd1 _09169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11200_ _11218_/A _11200_/B vssd1 vssd1 vccd1 vccd1 _16890_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_160_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _13461_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
X_11131_ hold5619/X _11789_/B _11130_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11131_/X
+ sky130_fd_sc_hd__o211a_1
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ hold5579/X _11156_/B _11061_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _11062_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3060 _14263_/X vssd1 vssd1 vccd1 vccd1 _17930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_289_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18018_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_216_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10013_ _16495_/Q _10013_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__and3_1
XFILLER_0_194_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3071 _17813_/Q vssd1 vssd1 vccd1 vccd1 hold3071/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3082 _17926_/Q vssd1 vssd1 vccd1 vccd1 hold3082/X sky130_fd_sc_hd__dlygate4sd3_1
X_15870_ _17741_/CLK _15870_/D vssd1 vssd1 vccd1 vccd1 _15870_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3093 _18113_/Q vssd1 vssd1 vccd1 vccd1 hold3093/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_218_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18201_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 _13971_/X vssd1 vssd1 vccd1 vccd1 _17790_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2381 _14691_/X vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14821_ hold1843/X _14828_/B _14820_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 _08263_/X vssd1 vssd1 vccd1 vccd1 _15766_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1680 _16226_/Q vssd1 vssd1 vccd1 vccd1 hold1680/X sky130_fd_sc_hd__dlygate4sd3_1
X_17540_ _18378_/CLK _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_1
X_14752_ _14984_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__or2_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1691 _15638_/Q vssd1 vssd1 vccd1 vccd1 hold1691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12231_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ hold2389/X _17688_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__mux2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ hold5625/X _11201_/B _10914_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10915_/X
+ sky130_fd_sc_hd__o211a_1
X_17471_ _17506_/CLK _17471_/D vssd1 vssd1 vccd1 vccd1 _17471_/Q sky130_fd_sc_hd__dfxtp_1
X_14683_ hold1731/X _14714_/B _14682_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _14683_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _13461_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16422_ _18389_/CLK _16422_/D vssd1 vssd1 vccd1 vccd1 _16422_/Q sky130_fd_sc_hd__dfxtp_1
X_13634_ hold2382/X _17665_/Q _13826_/C vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10846_ hold5479/X _11732_/B _10845_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _10846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16353_ _18296_/CLK _16353_/D vssd1 vssd1 vccd1 vccd1 _16353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ hold1536/X hold4285/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13566_/B sky130_fd_sc_hd__mux2_1
X_10777_ hold5178/X _11159_/B _10776_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _10777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15304_ _15304_/A _15304_/B vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12516_ _12960_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _17348_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16284_ _18237_/CLK _16284_/D vssd1 vssd1 vccd1 vccd1 _16284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13496_ hold1352/X hold4334/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13497_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ hold611/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__or2_1
X_18023_ _18055_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12447_ hold554/X _12445_/A _12445_/B _12446_/X _12436_/A vssd1 vssd1 vccd1 vccd1
+ hold81/A sky130_fd_sc_hd__o311a_1
XFILLER_0_129_1375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ hold903/X _15165_/B _15165_/Y _15050_/A vssd1 vssd1 vccd1 vccd1 hold904/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12378_ hold3683/X _13782_/A _12377_/X vssd1 vssd1 vccd1 vccd1 _12378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14117_ hold2550/X _14142_/B _14116_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11329_ hold4996/X _12308_/B _11328_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15097_ _15205_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14048_ _14782_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17807_ _17870_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15999_ _18404_/CLK _15999_/D vssd1 vssd1 vccd1 vccd1 hold842/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08540_ hold88/X hold128/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ _17738_/CLK _17738_/D vssd1 vssd1 vccd1 vccd1 _17738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ hold1687/X _08486_/B _08470_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _08471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17669_ _17701_/CLK _17669_/D vssd1 vssd1 vccd1 vccd1 _17669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _12424_/A hold777/X vssd1 vssd1 vccd1 vccd1 _16128_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5902 _16320_/Q vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5913 _18457_/Q vssd1 vssd1 vccd1 vccd1 hold5913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5924 _17542_/Q vssd1 vssd1 vccd1 vccd1 hold5924/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5935 _17544_/Q vssd1 vssd1 vccd1 vccd1 hold5935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold210 hold2/X vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__clkbuf_8
Xhold5946 _17556_/Q vssd1 vssd1 vccd1 vccd1 hold5946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 input22/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__buf_1
XFILLER_0_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5957 data_in[15] vssd1 vssd1 vccd1 vccd1 hold343/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5968 data_in[29] vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 la_data_in[17] vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold34/X vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5979 _18272_/Q vssd1 vssd1 vccd1 vccd1 hold5979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _14362_/A vssd1 vssd1 vccd1 vccd1 _12969_/A sky130_fd_sc_hd__buf_4
Xfanout712 _13037_/A vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__buf_2
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ hold4040/X _10010_/B _09924_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09925_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout723 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__buf_4
XFILLER_0_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_382_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout734 _09063_/A vssd1 vssd1 vccd1 vccd1 _09015_/A sky130_fd_sc_hd__clkbuf_4
Xfanout745 _08377_/A vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__buf_4
Xfanout756 _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__buf_4
X_09856_ hold4801/X _10049_/B _09855_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09856_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout767 _14538_/C1 vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_311_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout778 _08349_/A vssd1 vssd1 vccd1 vccd1 _13792_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_225_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 _13935_/A vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__buf_4
X_08807_ _09015_/A hold313/X vssd1 vssd1 vccd1 vccd1 _16022_/D sky130_fd_sc_hd__and2_1
XFILLER_0_225_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ hold4877/X _10601_/B _09786_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09787_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08738_ _12426_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _15989_/D sky130_fd_sc_hd__and2_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ hold215/X hold769/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__mux2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ hold3165/X hold4614/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ hold4433/X _12344_/B _11679_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11680_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10631_ _16701_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10631_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _13734_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ hold1923/X hold4195/X _11096_/S vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _12310_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _17257_/D sky130_fd_sc_hd__nor2_1
X_13281_ _13281_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__and2_1
XFILLER_0_84_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ hold874/X hold3797/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15020_ hold331/X hold393/X vssd1 vssd1 vccd1 vccd1 hold394/A sky130_fd_sc_hd__or2_1
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12232_ hold4281/X _12347_/B _12231_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12163_ hold5455/X _12353_/B _12162_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ hold2244/X _16862_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__mux2_1
X_12094_ hold5413/X _12353_/B _12093_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _12094_/X
+ sky130_fd_sc_hd__o211a_1
X_16971_ _18425_/CLK _16971_/D vssd1 vssd1 vccd1 vccd1 _16971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _17286_/CLK _15922_/D vssd1 vssd1 vccd1 vccd1 hold676/A sky130_fd_sc_hd__dfxtp_1
X_11045_ hold2581/X _16839_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _17712_/CLK _15853_/D vssd1 vssd1 vccd1 vccd1 _15853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14804_ _15197_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15784_ _17737_/CLK _15784_/D vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12996_ _12996_/A _12996_/B vssd1 vssd1 vccd1 vccd1 _17508_/D sky130_fd_sc_hd__and2_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17523_ _17523_/CLK hold959/X vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_235_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ _14735_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14784_/B sky130_fd_sc_hd__or2_4
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ hold4145/X _13871_/B _11946_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _14774_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14666_/Y sky130_fd_sc_hd__nand2_1
X_17454_ _17455_/CLK _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11878_ hold5443/X _13862_/B _11877_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _11878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16405_ _18316_/CLK _16405_/D vssd1 vssd1 vccd1 vccd1 _16405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13617_ _13800_/A _13617_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10829_ hold1666/X _16767_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14597_ hold2484/X _14612_/B _14596_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14597_/X
+ sky130_fd_sc_hd__o211a_1
X_17385_ _18434_/CLK _17385_/D vssd1 vssd1 vccd1 vccd1 _17385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ _18389_/CLK _16336_/D vssd1 vssd1 vccd1 vccd1 _16336_/Q sky130_fd_sc_hd__dfxtp_1
X_13548_ _13761_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16267_ _17499_/CLK _16267_/D vssd1 vssd1 vccd1 vccd1 _16267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _13734_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5209 _11269_/X vssd1 vssd1 vccd1 vccd1 _16913_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15218_ hold964/X _15221_/B _15217_/Y _15058_/A vssd1 vssd1 vccd1 vccd1 hold965/A
+ sky130_fd_sc_hd__o211a_1
X_18006_ _18006_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _17479_/CLK _16198_/D vssd1 vssd1 vccd1 vccd1 _16198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4508 _13777_/X vssd1 vssd1 vccd1 vccd1 _17712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4519 _17151_/Q vssd1 vssd1 vccd1 vccd1 hold4519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15203_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3807 _10864_/X vssd1 vssd1 vccd1 vccd1 _16778_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3818 _10303_/X vssd1 vssd1 vccd1 vccd1 _16591_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3829 _16932_/Q vssd1 vssd1 vccd1 vccd1 hold3829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07971_ hold2548/X _07978_/B _07970_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _07971_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_226_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09710_ _18305_/Q _16394_/Q _11159_/C vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09641_ hold3015/X _16371_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_235_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09572_ hold986/X _13254_/A _10190_/S vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _08730_/A _13046_/C vssd1 vssd1 vccd1 vccd1 _08528_/S sky130_fd_sc_hd__or2_2
XFILLER_0_195_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _15513_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _15824_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09006_ hold113/X hold281/X _09006_/S vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__mux2_1
Xhold5710 _13627_/X vssd1 vssd1 vccd1 vccd1 _17662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5721 _17634_/Q vssd1 vssd1 vccd1 vccd1 hold5721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5732 _13546_/X vssd1 vssd1 vccd1 vccd1 _17635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5743 _17600_/Q vssd1 vssd1 vccd1 vccd1 hold5743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5754 _13348_/X vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5765 hold5923/X vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5776 output85/X vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5787 hold5939/X vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5798 output84/X vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_40_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 _09340_/X vssd1 vssd1 vccd1 vccd1 _15490_/B1 sky130_fd_sc_hd__buf_8
Xfanout531 _09177_/A2 vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout542 _08448_/Y vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__buf_8
X_09908_ hold2997/X hold3898/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_217_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout553 _08228_/Y vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__buf_8
XFILLER_0_233_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout564 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__clkbuf_8
Xfanout575 _14610_/B vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__buf_6
Xfanout586 _13225_/B vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__buf_4
X_09839_ _18348_/Q hold3858/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__mux2_1
Xfanout597 _12985_/S vssd1 vssd1 vccd1 vccd1 _12997_/S sky130_fd_sc_hd__buf_6
XFILLER_0_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12850_ hold1227/X hold3304/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_214_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _17091_/Q _11801_/B _12365_/C vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__and3_1
XFILLER_0_197_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ hold2063/X hold3308/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__mux2_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ hold3120/X _14541_/B _14519_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14520_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ hold915/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14451_/X sky130_fd_sc_hd__or2_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11663_ hold1973/X _17045_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13402_ hold4334/X _13880_/B _13401_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13402_/X
+ sky130_fd_sc_hd__o211a_1
X_10614_ hold3549/X _10536_/A _10613_/X vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17170_ _17170_/CLK _17170_/D vssd1 vssd1 vccd1 vccd1 _17170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14382_ _15072_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ hold2463/X _17022_/Q _11594_/S vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__mux2_1
X_16121_ _17340_/CLK _16121_/D vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13333_ hold5080/X _13811_/B _13332_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10545_ _10998_/A _10545_/B vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16052_ _17330_/CLK _16052_/D vssd1 vssd1 vccd1 vccd1 hold443/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13264_ _13257_/X _13263_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_228_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10476_ _10476_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ hold966/X hold514/X _15002_/Y _15058_/A vssd1 vssd1 vccd1 vccd1 hold967/A
+ sky130_fd_sc_hd__o211a_1
X_12215_ hold1585/X _17229_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _12216_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13195_ _13194_/X _16917_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_233_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18193_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ hold2586/X hold5599/X _12338_/C vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12077_ hold2164/X _17183_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__mux2_1
X_16954_ _17896_/CLK _16954_/D vssd1 vssd1 vccd1 vccd1 _16954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15905_ _16095_/CLK _15905_/D vssd1 vssd1 vccd1 vccd1 hold438/A sky130_fd_sc_hd__dfxtp_1
X_11028_ _11124_/A _11028_/B vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__or2_1
X_16885_ _18054_/CLK _16885_/D vssd1 vssd1 vccd1 vccd1 _16885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _17729_/CLK _15836_/D vssd1 vssd1 vccd1 vccd1 _15836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _17726_/CLK _15767_/D vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfxtp_1
X_12979_ hold2630/X hold3138/X _12985_/S vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__mux2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ _17506_/CLK _17506_/D vssd1 vssd1 vccd1 vccd1 _17506_/Q sky130_fd_sc_hd__dfxtp_1
X_14718_ _15004_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15698_ _17266_/CLK _15698_/D vssd1 vssd1 vccd1 vccd1 _15698_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _18436_/CLK _17437_/D vssd1 vssd1 vccd1 vccd1 _17437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14649_ hold3097/X _14664_/B _14648_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14649_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_16 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_27 _08963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08170_ _15521_/A hold2074/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__mux2_1
XANTENNA_38 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _17370_/CLK _17368_/D vssd1 vssd1 vccd1 vccd1 _17368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_49 _15555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16319_ _16320_/CLK _16319_/D vssd1 vssd1 vccd1 vccd1 _16319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17299_ _17299_/CLK _17299_/D vssd1 vssd1 vccd1 vccd1 hold795/A sky130_fd_sc_hd__dfxtp_1
Xhold5006 _17258_/Q vssd1 vssd1 vccd1 vccd1 hold5006/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5017 _10699_/X vssd1 vssd1 vccd1 vccd1 _16723_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5028 _16964_/Q vssd1 vssd1 vccd1 vccd1 hold5028/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput101 _13113_/A vssd1 vssd1 vccd1 vccd1 hold5806/A sky130_fd_sc_hd__buf_6
Xhold5039 _09754_/X vssd1 vssd1 vccd1 vccd1 _16408_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4305 _17233_/Q vssd1 vssd1 vccd1 vccd1 hold4305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput112 hold5848/X vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_12
Xhold4316 _13564_/X vssd1 vssd1 vccd1 vccd1 _17641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput123 hold5892/X vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_12
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput134 hold5867/X vssd1 vssd1 vccd1 vccd1 hold5868/A sky130_fd_sc_hd__buf_6
Xhold4327 _17089_/Q vssd1 vssd1 vccd1 vccd1 hold4327/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput145 hold5859/X vssd1 vssd1 vccd1 vccd1 hold5860/A sky130_fd_sc_hd__buf_6
Xhold4338 _17605_/Q vssd1 vssd1 vccd1 vccd1 hold4338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3604 _16720_/Q vssd1 vssd1 vccd1 vccd1 hold3604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4349 _13459_/X vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3615 _16333_/Q vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3626 _12360_/Y vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3637 _17578_/Q vssd1 vssd1 vccd1 vccd1 hold3637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3648 _13857_/Y vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2903 _17845_/Q vssd1 vssd1 vccd1 vccd1 hold2903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3659 _16553_/Q vssd1 vssd1 vccd1 vccd1 hold3659/X sky130_fd_sc_hd__buf_1
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2914 _15556_/X vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2925 _17794_/Q vssd1 vssd1 vccd1 vccd1 hold2925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2936 _14815_/X vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07954_ _14517_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2947 _18397_/Q vssd1 vssd1 vccd1 vccd1 hold2947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2958 _14301_/X vssd1 vssd1 vccd1 vccd1 _17948_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2969 _15571_/Q vssd1 vssd1 vccd1 vccd1 hold2969/X sky130_fd_sc_hd__dlygate4sd3_1
X_07885_ hold202/X _14789_/A vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__or2_4
XFILLER_0_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _09984_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_29_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_29_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _09963_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_214_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08506_ hold1320/X _08503_/Y _08505_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08506_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09486_ hold1833/X _09483_/X _09485_/Y vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08437_ _14330_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _15537_/A hold2379/X hold134/X vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08299_ _14517_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ hold5236/X _11095_/A2 _10329_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_239_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5540 _10828_/X vssd1 vssd1 vccd1 vccd1 _16766_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10261_ hold3874/X _10646_/B _10260_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5551 _16848_/Q vssd1 vssd1 vccd1 vccd1 hold5551/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5562 _11377_/X vssd1 vssd1 vccd1 vccd1 _16949_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5573 _16771_/Q vssd1 vssd1 vccd1 vccd1 hold5573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5584 _11041_/X vssd1 vssd1 vccd1 vccd1 _16837_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12000_ _13797_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__or2_1
Xhold4850 _10408_/X vssd1 vssd1 vccd1 vccd1 _16626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5595 _17055_/Q vssd1 vssd1 vccd1 vccd1 hold5595/X sky130_fd_sc_hd__dlygate4sd3_1
X_10192_ hold5665/X _10070_/B _10191_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10192_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4861 _16857_/Q vssd1 vssd1 vccd1 vccd1 hold4861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4872 _12324_/Y vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4883 _16508_/Q vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4894 _11101_/X vssd1 vssd1 vccd1 vccd1 _16857_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout350 _08759_/S vssd1 vssd1 vccd1 vccd1 _08793_/S sky130_fd_sc_hd__buf_8
XFILLER_0_22_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout361 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15221_/B sky130_fd_sc_hd__buf_8
XFILLER_0_205_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout372 hold513/X vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__clkbuf_1
Xfanout383 _14784_/B vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__buf_8
X_13951_ hold1119/X _13995_/A2 _13950_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _13951_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout394 _14501_/Y vssd1 vssd1 vccd1 vccd1 _14535_/B sky130_fd_sc_hd__buf_8
X_12902_ hold3167/X _12901_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__mux2_1
X_16670_ _18226_/CLK _16670_/D vssd1 vssd1 vccd1 vccd1 _16670_/Q sky130_fd_sc_hd__dfxtp_1
X_13882_ _13888_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _17747_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15621_ _17217_/CLK _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ hold3367/X _12832_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18340_ _18380_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12764_ hold3815/X _12763_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__mux2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ hold1292/X _15560_/A2 _15551_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _15552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14968_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11715_ _12213_/A _11715_/B vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__or2_1
X_15483_ hold790/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18271_ _18303_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ hold3785/X _12694_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__mux2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _17623_/CLK _17222_/D vssd1 vssd1 vccd1 vccd1 _17222_/Q sky130_fd_sc_hd__dfxtp_1
X_14434_ hold2705/X _14433_/B _14433_/Y _14434_/C1 vssd1 vssd1 vccd1 vccd1 _14434_/X
+ sky130_fd_sc_hd__o211a_1
X_11646_ _11652_/A _11646_/B vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 input14/A vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_0_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 input25/A vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_6
X_14365_ _15099_/A hold2978/X hold333/X vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__mux2_1
X_17153_ _17153_/CLK _17153_/D vssd1 vssd1 vccd1 vccd1 _17153_/Q sky130_fd_sc_hd__dfxtp_1
Xinput36 input36/A vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11577_ _11679_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_414_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17842_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 input47/A vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
X_16104_ _17327_/CLK _16104_/D vssd1 vssd1 vccd1 vccd1 hold480/A sky130_fd_sc_hd__dfxtp_1
Xinput58 input58/A vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_6
X_13316_ hold1088/X hold3890/X _13412_/S vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput69 input69/A vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
X_10528_ hold3766/X _10622_/B _10527_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10528_/X
+ sky130_fd_sc_hd__o211a_1
X_17084_ _17265_/CLK _17084_/D vssd1 vssd1 vccd1 vccd1 _17084_/Q sky130_fd_sc_hd__dfxtp_1
X_14296_ hold926/X _14336_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__or2_1
Xhold809 hold809/A vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _13311_/A1 _13245_/X _13246_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13247_/X
+ sky130_fd_sc_hd__o211a_1
X_16035_ _17299_/CLK _16035_/D vssd1 vssd1 vccd1 vccd1 hold610/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10459_ hold3776/X _10477_/A2 _10458_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13178_ _17573_/Q _17107_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12129_ _13797_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or2_1
X_17986_ _18018_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 hold426/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1509 _18129_/Q vssd1 vssd1 vccd1 vccd1 hold1509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16937_ _17815_/CLK _16937_/D vssd1 vssd1 vccd1 vccd1 _16937_/Q sky130_fd_sc_hd__dfxtp_1
X_16868_ _18071_/CLK _16868_/D vssd1 vssd1 vccd1 vccd1 _16868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ _17425_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 _15819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16799_ _18067_/CLK _16799_/D vssd1 vssd1 vccd1 vccd1 _16799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _18458_/Q _07802_/B _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09271_ hold367/X _16247_/Q _09273_/S vssd1 vssd1 vccd1 vccd1 hold535/A sky130_fd_sc_hd__mux2_1
XFILLER_0_158_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08222_ hold2772/X _08209_/B _08221_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _08222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17306_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _14878_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4102 _13417_/X vssd1 vssd1 vccd1 vccd1 _17592_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4113 _15463_/X vssd1 vssd1 vccd1 vccd1 _15464_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4124 _09598_/X vssd1 vssd1 vccd1 vccd1 _16356_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4135 _17671_/Q vssd1 vssd1 vccd1 vccd1 hold4135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4146 _11947_/X vssd1 vssd1 vccd1 vccd1 _17139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3401 _16874_/Q vssd1 vssd1 vccd1 vccd1 hold3401/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3412 _16391_/Q vssd1 vssd1 vccd1 vccd1 hold3412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4157 _17390_/Q vssd1 vssd1 vccd1 vccd1 hold4157/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3423 _09523_/X vssd1 vssd1 vccd1 vccd1 _16331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4168 _17405_/Q vssd1 vssd1 vccd1 vccd1 hold4168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3434 _17181_/Q vssd1 vssd1 vccd1 vccd1 hold3434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4179 _17003_/Q vssd1 vssd1 vccd1 vccd1 hold4179/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3445 _10948_/X vssd1 vssd1 vccd1 vccd1 _16806_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2700 _08402_/X vssd1 vssd1 vccd1 vccd1 _15831_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3456 _17178_/Q vssd1 vssd1 vccd1 vccd1 hold3456/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2711 _17797_/Q vssd1 vssd1 vccd1 vccd1 hold2711/X sky130_fd_sc_hd__dlygate4sd3_1
X_08986_ _12436_/A hold349/X vssd1 vssd1 vccd1 vccd1 _16110_/D sky130_fd_sc_hd__and2_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2722 _14460_/X vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3467 _12659_/X vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2733 _18026_/Q vssd1 vssd1 vccd1 vccd1 hold2733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3478 _17216_/Q vssd1 vssd1 vccd1 vccd1 hold3478/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3489 _12569_/X vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2744 _07965_/X vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2755 _18335_/Q vssd1 vssd1 vccd1 vccd1 hold2755/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ hold1746/X _07924_/B _07936_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _07937_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2766 _18369_/Q vssd1 vssd1 vccd1 vccd1 hold2766/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2777 _14101_/X vssd1 vssd1 vccd1 vccd1 _17853_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2788 _14679_/X vssd1 vssd1 vccd1 vccd1 _18130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 _18304_/Q vssd1 vssd1 vccd1 vccd1 hold2799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07868_ hold2890/X _07869_/B _07867_/Y _08149_/A vssd1 vssd1 vccd1 vccd1 _07868_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09607_ hold3412/X _10025_/B _09606_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07799_ _11158_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_195_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ hold5052/X _10034_/B _09537_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _09472_/B _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__and3_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ hold5507/X _12329_/B _11499_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _11500_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _17333_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ hold4990/X _12299_/B _11430_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11431_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _15549_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ hold5352/X _11732_/B _11361_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11362_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _13100_/X hold4616/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__mux2_1
X_10313_ hold2365/X hold3944/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14081_ hold2985/X _14094_/B _14080_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ hold4364/X _12338_/B _11292_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11293_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13032_ _13056_/C hold922/X hold958/A vssd1 vssd1 vccd1 vccd1 _13032_/Y sky130_fd_sc_hd__o21ai_1
Xhold5370 _17558_/Q vssd1 vssd1 vccd1 vccd1 hold5370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5381 _16601_/Q vssd1 vssd1 vccd1 vccd1 hold5381/X sky130_fd_sc_hd__dlygate4sd3_1
X_10244_ hold2341/X _16572_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5392 _11836_/X vssd1 vssd1 vccd1 vccd1 _17102_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4680 _11721_/Y vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17840_ _17862_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10175_ hold1813/X hold4775/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__mux2_1
Xhold4691 _17103_/Q vssd1 vssd1 vccd1 vccd1 hold4691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3990 _16663_/Q vssd1 vssd1 vccd1 vccd1 hold3990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17771_ _17890_/CLK hold126/X vssd1 vssd1 vccd1 vccd1 _17771_/Q sky130_fd_sc_hd__dfxtp_1
X_14983_ hold1283/X hold514/X _14982_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14983_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout180 _11168_/B vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout191 _13886_/B vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16722_ _18018_/CLK _16722_/D vssd1 vssd1 vccd1 vccd1 _16722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13934_ _14328_/A hold2060/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13935_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16653_ _18209_/CLK _16653_/D vssd1 vssd1 vccd1 vccd1 _16653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _17742_/Q _13871_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _17897_/CLK _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12816_ _12912_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _17448_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16584_ _18263_/CLK _16584_/D vssd1 vssd1 vccd1 vccd1 _16584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ hold1434/X _17719_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ _18323_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _15535_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _17425_/D sky130_fd_sc_hd__and2_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18254_ _18382_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15466_ hold456/X _09386_/A _09386_/D _15904_/Q vssd1 vssd1 vccd1 vccd1 _15471_/B
+ sky130_fd_sc_hd__a22o_1
X_12678_ _12810_/A _12678_/B vssd1 vssd1 vccd1 vccd1 _17402_/D sky130_fd_sc_hd__and2_1
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17205_ _17269_/CLK _17205_/D vssd1 vssd1 vccd1 vccd1 _17205_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ hold4014/X _11726_/B _11628_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11629_/X
+ sky130_fd_sc_hd__o211a_1
X_14417_ _15205_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__or2_1
X_18185_ _18199_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15397_ hold186/X _09357_/A _09386_/D hold618/X _15396_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17136_ _17718_/CLK _17136_/D vssd1 vssd1 vccd1 vccd1 _17136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14348_ _14348_/A _14348_/B vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__and2_1
Xhold606 input19/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold617 hold617/A vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold628 hold628/A vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold639 hold639/A vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17067_ _18425_/CLK _17067_/D vssd1 vssd1 vccd1 vccd1 _17067_/Q sky130_fd_sc_hd__dfxtp_1
X_14279_ hold2759/X _14272_/B _14278_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16018_ _17335_/CLK _16018_/D vssd1 vssd1 vccd1 vccd1 hold563/A sky130_fd_sc_hd__dfxtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _14566_/X vssd1 vssd1 vccd1 vccd1 hold2007/X sky130_fd_sc_hd__dlygate4sd3_1
X_08840_ hold568/X hold878/X _08866_/S vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__mux2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 _08030_/X vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _15858_/Q vssd1 vssd1 vccd1 vccd1 hold2029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _08178_/X vssd1 vssd1 vccd1 vccd1 _15725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08771_ hold353/X hold484/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__mux2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _08118_/X vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1328 _09290_/X vssd1 vssd1 vccd1 vccd1 _16255_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _18064_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1339 _14739_/X vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09323_ _15219_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_336_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09254_ _12738_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _16238_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08205_ _15539_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08205_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ hold2562/X _09218_/B _09184_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _09185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ hold469/X hold590/X hold240/X vssd1 vssd1 vccd1 vccd1 hold591/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08067_ hold2592/X _08097_/A2 _08066_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3220 _18029_/Q vssd1 vssd1 vccd1 vccd1 hold3220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3231 _12593_/X vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3242 _16331_/Q vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3253 _17494_/Q vssd1 vssd1 vccd1 vccd1 hold3253/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3264 _17486_/Q vssd1 vssd1 vccd1 vccd1 hold3264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2530 _14041_/X vssd1 vssd1 vccd1 vccd1 _17824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3275 _17373_/Q vssd1 vssd1 vccd1 vccd1 hold3275/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3286 _17377_/Q vssd1 vssd1 vccd1 vccd1 hold3286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2541 _14147_/X vssd1 vssd1 vccd1 vccd1 _17875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2552 _15702_/Q vssd1 vssd1 vccd1 vccd1 hold2552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3297 _17464_/Q vssd1 vssd1 vccd1 vccd1 hold3297/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17822_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08969_ hold379/X hold678/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__mux2_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 _09185_/X vssd1 vssd1 vccd1 vccd1 _16204_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2574 _14047_/X vssd1 vssd1 vccd1 vccd1 _17827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1840 _14817_/X vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2585 _16238_/Q vssd1 vssd1 vccd1 vccd1 hold2585/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1851 _18386_/Q vssd1 vssd1 vccd1 vccd1 hold1851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2596 _15812_/Q vssd1 vssd1 vccd1 vccd1 hold2596/X sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ hold4071/X _13871_/B _11979_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11980_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1862 _14159_/X vssd1 vssd1 vccd1 vccd1 _17881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 _17793_/Q vssd1 vssd1 vccd1 vccd1 hold1873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1884 _14293_/X vssd1 vssd1 vccd1 vccd1 _17944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1895 _17911_/Q vssd1 vssd1 vccd1 vccd1 hold1895/X sky130_fd_sc_hd__dlygate4sd3_1
X_10931_ hold3112/X hold4523/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ hold1056/X _16778_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__mux2_1
X_13650_ _13746_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13650_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ hold1296/X _17378_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__mux2_1
X_13581_ _13776_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ hold3110/X hold5016/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__mux2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ hold158/X _15486_/A2 _09357_/B _16061_/Q vssd1 vssd1 vccd1 vccd1 _15320_/X
+ sky130_fd_sc_hd__a22o_1
X_12532_ hold2535/X hold3274/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12463_ hold26/X _12445_/A _12445_/B _12462_/X _15324_/A vssd1 vssd1 vccd1 vccd1
+ hold27/A sky130_fd_sc_hd__o311a_1
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _16289_/Q _15477_/A2 _15487_/B1 hold627/X _15250_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11414_ hold2697/X hold3525/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__mux2_1
X_14202_ _14774_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__nand2_1
X_15182_ _15182_/A hold393/X vssd1 vssd1 vccd1 vccd1 _15211_/B sky130_fd_sc_hd__or2_4
X_12394_ _15264_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _17290_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ hold2463/X _14148_/B _14132_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _14133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ hold2331/X hold4069/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _14403_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11276_ hold2155/X hold4793/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11277_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_219_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _15519_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__or2_1
X_10227_ _10497_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__or2_1
XTAP_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _17855_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10158_ _10536_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17754_ _18017_/CLK _17754_/D vssd1 vssd1 vccd1 vccd1 _17754_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _10563_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__or2_1
X_14966_ hold754/X hold393/X vssd1 vssd1 vccd1 vccd1 hold513/A sky130_fd_sc_hd__nor2_1
XFILLER_0_234_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16705_ _18229_/CLK _16705_/D vssd1 vssd1 vccd1 vccd1 _16705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ _13917_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _17764_/D sky130_fd_sc_hd__and2_1
X_17685_ _17749_/CLK _17685_/D vssd1 vssd1 vccd1 vccd1 _17685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14897_ _14897_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__or2_2
XFILLER_0_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ _18180_/CLK _16636_/D vssd1 vssd1 vccd1 vccd1 _16636_/Q sky130_fd_sc_hd__dfxtp_1
X_13848_ hold3306/X _13746_/A _13847_/X vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16567_ _16631_/CLK _16567_/D vssd1 vssd1 vccd1 vccd1 _16567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13779_ _13779_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ _18370_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15518_ hold2081/X _15507_/Y _15517_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _15518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16498_ _18377_/CLK _16498_/D vssd1 vssd1 vccd1 vccd1 _16498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18237_ _18237_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15449_ hold127/X _15484_/A2 _15447_/X vssd1 vssd1 vccd1 vccd1 _15452_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_143_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _18232_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17903_/CLK _17119_/D vssd1 vssd1 vccd1 vccd1 _17119_/Q sky130_fd_sc_hd__dfxtp_1
Xhold425 hold425/A vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _18131_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
Xhold436 hold436/A vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold447 hold447/A vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09941_ hold1648/X hold4739/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09942_/B sky130_fd_sc_hd__mux2_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout905 hold719/X vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__buf_12
Xfanout916 hold559/X vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__clkbuf_16
Xfanout927 _15213_/A vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__buf_12
XFILLER_0_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09872_ hold1885/X hold4765/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 hold1248/X vssd1 vssd1 vccd1 vccd1 hold1249/A sky130_fd_sc_hd__buf_6
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08823_ _12386_/A hold301/X vssd1 vssd1 vccd1 vccd1 _16030_/D sky130_fd_sc_hd__and2_1
Xhold1103 _15114_/X vssd1 vssd1 vccd1 vccd1 _18339_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 _09069_/X vssd1 vssd1 vccd1 vccd1 _16149_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _18440_/Q vssd1 vssd1 vccd1 vccd1 hold1125/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1136 input43/X vssd1 vssd1 vccd1 vccd1 hold1136/X sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _15414_/A hold362/X vssd1 vssd1 vccd1 vccd1 _15997_/D sky130_fd_sc_hd__and2_1
Xhold1147 _18220_/Q vssd1 vssd1 vccd1 vccd1 hold1147/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1158 _09123_/X vssd1 vssd1 vccd1 vccd1 _16175_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1169 _15001_/X vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08685_ hold98/X hold781/X _08685_/S vssd1 vssd1 vccd1 vccd1 hold782/A sky130_fd_sc_hd__mux2_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_170_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18060_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09306_ hold1090/X _09325_/B _09305_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ _15513_/A hold2745/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09168_ _15551_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08119_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ hold2894/X _09106_/B _09098_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _09099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_222_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11130_ _11670_/A _11130_/B vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__or2_1
Xhold970 hold977/X vssd1 vssd1 vccd1 vccd1 hold978/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3050 _09197_/X vssd1 vssd1 vccd1 vccd1 _16210_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ _11203_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _16494_/D sky130_fd_sc_hd__nor2_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3061 _17787_/Q vssd1 vssd1 vccd1 vccd1 hold3061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3072 _14019_/X vssd1 vssd1 vccd1 vccd1 _17813_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3083 _14255_/X vssd1 vssd1 vccd1 vccd1 _17926_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3094 _14645_/X vssd1 vssd1 vccd1 vccd1 _18113_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2360 _08216_/X vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _15213_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__or2_1
Xhold2371 _18102_/Q vssd1 vssd1 vccd1 vccd1 hold2371/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 _15798_/Q vssd1 vssd1 vccd1 vccd1 hold2382/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2393 _16165_/Q vssd1 vssd1 vccd1 vccd1 hold2393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 _15586_/Q vssd1 vssd1 vccd1 vccd1 hold1670/X sky130_fd_sc_hd__dlygate4sd3_1
X_14751_ hold1945/X _14774_/B _14750_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14751_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1681 _09229_/X vssd1 vssd1 vccd1 vccd1 _16226_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1692 _07991_/X vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11963_ hold2210/X hold4125/X _13868_/C vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_258_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18065_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ hold4089/X _13814_/B _13701_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _13702_/X
+ sky130_fd_sc_hd__o211a_1
X_10914_ _11106_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__or2_1
X_17470_ _17506_/CLK _17470_/D vssd1 vssd1 vccd1 vccd1 _17470_/Q sky130_fd_sc_hd__dfxtp_1
X_14682_ _14968_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14682_/X sky130_fd_sc_hd__or2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ hold2117/X hold3639/X _13556_/S vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _18364_/CLK _16421_/D vssd1 vssd1 vccd1 vccd1 _16421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13633_ hold5755/X _13832_/B _13632_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13633_/X
+ sky130_fd_sc_hd__o211a_1
X_10845_ _11553_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _18108_/CLK _16352_/D vssd1 vssd1 vccd1 vccd1 _16352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10776_ _11064_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__or2_1
X_13564_ hold4315/X _13880_/B _13563_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13564_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _15490_/A1 _15295_/X _15302_/X _15490_/B1 hold5832/A vssd1 vssd1 vccd1 vccd1
+ _15303_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12515_ _07826_/A _12514_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16283_ _18459_/CLK _16283_/D vssd1 vssd1 vccd1 vccd1 _16283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13495_ hold4303/X _13880_/B _13494_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ _18054_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12446_ _17316_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__or2_1
X_15234_ hold2947/X _15221_/B _15233_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15234_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15165_ _15219_/A _15165_/B vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__nand2_1
X_12377_ _17283_/Q _13877_/B _13877_/C vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__and3_1
XFILLER_0_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11328_ _12213_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__or2_1
X_14116_ _14116_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__or2_1
X_15096_ hold1660/X _15111_/B _15095_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15096_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14047_ hold2573/X _14038_/B _14046_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _14047_/X
+ sky130_fd_sc_hd__o211a_1
X_11259_ _11643_/A _11259_/B vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _17891_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _18411_/CLK _15998_/D vssd1 vssd1 vccd1 vccd1 _15998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _17737_/CLK _17737_/D vssd1 vssd1 vccd1 vccd1 _17737_/Q sky130_fd_sc_hd__dfxtp_1
X_14949_ hold986/X _14952_/B _14948_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 hold987/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08470_ _15203_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08470_/X sky130_fd_sc_hd__or2_1
X_17668_ _17700_/CLK _17668_/D vssd1 vssd1 vccd1 vccd1 _17668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16619_ _18175_/CLK _16619_/D vssd1 vssd1 vccd1 vccd1 _16619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17599_ _17729_/CLK _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09022_ hold361/X hold776/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold777/A sky130_fd_sc_hd__mux2_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5903 _09477_/X vssd1 vssd1 vccd1 vccd1 _09483_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5914 _07793_/X vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold200 hold530/X vssd1 vssd1 vccd1 vccd1 hold531/A sky130_fd_sc_hd__buf_4
Xhold5925 _17548_/Q vssd1 vssd1 vccd1 vccd1 hold5925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5936 _17543_/Q vssd1 vssd1 vccd1 vccd1 hold5936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5947 _17528_/Q vssd1 vssd1 vccd1 vccd1 hold5947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold14/X vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__buf_4
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5958 data_in[25] vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 input45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5969 becStatus[1] vssd1 vssd1 vccd1 vccd1 hold951/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 input12/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__buf_1
XFILLER_0_106_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _09933_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__or2_1
Xfanout702 _14362_/A vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__buf_4
Xfanout713 _13037_/A vssd1 vssd1 vccd1 vccd1 _12436_/A sky130_fd_sc_hd__buf_4
Xfanout724 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _12404_/A sky130_fd_sc_hd__buf_2
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout735 _09063_/A vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__buf_2
XFILLER_0_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout746 _08377_/A vssd1 vssd1 vccd1 vccd1 _13483_/C1 sky130_fd_sc_hd__buf_2
X_09855_ _09954_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__or2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 fanout770/X vssd1 vssd1 vccd1 vccd1 _12073_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _14538_/C1 vssd1 vssd1 vccd1 vccd1 _14472_/C1 sky130_fd_sc_hd__buf_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 fanout796/X vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ hold312/X _16022_/Q _08866_/S vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__mux2_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _10488_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__or2_1
XFILLER_0_225_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ hold113/X hold767/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__mux2_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_351_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17642_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08668_ _12418_/A hold414/X vssd1 vssd1 vccd1 vccd1 _15955_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ hold554/X hold676/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold677/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ _11218_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _16700_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ hold4795/X _10571_/B _10560_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _10561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ hold4672/X _12204_/A _12299_/X vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13280_ _13273_/X _13279_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10492_ hold5262/X _10625_/B _10491_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _12231_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ _13794_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ hold5553/X _11207_/B _11112_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12093_ _13794_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__or2_1
X_16970_ _17816_/CLK _16970_/D vssd1 vssd1 vccd1 vccd1 _16970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15921_ _18406_/CLK _15921_/D vssd1 vssd1 vccd1 vccd1 hold582/A sky130_fd_sc_hd__dfxtp_1
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11044_ hold4219/X _11729_/B _11043_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _11044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_439_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _17647_/CLK _15852_/D vssd1 vssd1 vccd1 vccd1 _15852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _17959_/Q vssd1 vssd1 vccd1 vccd1 hold2190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14803_ hold1161/X _14826_/B _14802_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14803_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _17650_/CLK _15783_/D vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ hold3254/X _12994_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__mux2_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17523_/CLK _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14734_ _14735_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nor2_2
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _12267_/A _11946_/B vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__or2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17455_/CLK _17453_/D vssd1 vssd1 vccd1 vccd1 _17453_/Q sky130_fd_sc_hd__dfxtp_1
X_14665_ hold1954/X _14664_/B _14664_/Y _14815_/C1 vssd1 vssd1 vccd1 vccd1 _14665_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _12261_/A _11877_/B vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__or2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16404_ _18321_/CLK _16404_/D vssd1 vssd1 vccd1 vccd1 _16404_/Q sky130_fd_sc_hd__dfxtp_1
X_13616_ hold2315/X _17659_/Q _13622_/S vssd1 vssd1 vccd1 vccd1 _13617_/B sky130_fd_sc_hd__mux2_1
X_17384_ _18434_/CLK _17384_/D vssd1 vssd1 vccd1 vccd1 _17384_/Q sky130_fd_sc_hd__dfxtp_1
X_10828_ hold5539/X _11762_/B _10827_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _10828_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14596_ _14758_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14596_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ _18366_/CLK _16335_/D vssd1 vssd1 vccd1 vccd1 _16335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13547_ hold663/X hold4545/X _13856_/C vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10759_ hold4336/X _11147_/B _10758_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ _17370_/CLK _16266_/D vssd1 vssd1 vccd1 vccd1 _16266_/Q sky130_fd_sc_hd__dfxtp_1
X_13478_ hold2482/X _17613_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__mux2_1
X_18005_ _18071_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
X_15217_ _15217_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12429_ hold578/X hold620/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16197_ _17481_/CLK _16197_/D vssd1 vssd1 vccd1 vccd1 _16197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4509 _16765_/Q vssd1 vssd1 vccd1 vccd1 hold4509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15148_ hold3134/X _15167_/B _15147_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _15148_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3808 _16364_/Q vssd1 vssd1 vccd1 vccd1 hold3808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3819 _16476_/Q vssd1 vssd1 vccd1 vccd1 hold3819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_239_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07970_ _15539_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__or2_1
X_15079_ hold746/X _15125_/B vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09640_ hold5621/X _11201_/B _09639_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09640_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18403_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09571_ hold3653/X _10049_/B _09570_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09571_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_19_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_19_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08522_ hold990/X _13043_/C vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_223_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ hold1061/X _08488_/B _08452_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08384_ _14726_/A hold2264/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09005_ _09061_/A hold216/X vssd1 vssd1 vccd1 vccd1 _16119_/D sky130_fd_sc_hd__and2_1
Xhold5700 _09976_/X vssd1 vssd1 vccd1 vccd1 _16482_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5711 _16554_/Q vssd1 vssd1 vccd1 vccd1 hold5711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5722 _13447_/X vssd1 vssd1 vccd1 vccd1 _17602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5733 _17678_/Q vssd1 vssd1 vccd1 vccd1 hold5733/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5744 _13345_/X vssd1 vssd1 vccd1 vccd1 _17568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5755 _17696_/Q vssd1 vssd1 vccd1 vccd1 hold5755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5766 output74/X vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_12
Xhold5777 hold5930/X vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5788 output92/X vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_12
Xhold5799 hold5935/X vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout510 _10481_/S vssd1 vssd1 vccd1 vccd1 _10601_/C sky130_fd_sc_hd__clkbuf_8
Xclkbuf_6_58_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_58_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xfanout521 _09340_/X vssd1 vssd1 vccd1 vccd1 _15481_/B1 sky130_fd_sc_hd__clkbuf_4
X_09907_ hold3868/X _10025_/B _09906_/X _14915_/C1 vssd1 vssd1 vccd1 vccd1 _09907_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout532 _09124_/Y vssd1 vssd1 vccd1 vccd1 _09177_/A2 sky130_fd_sc_hd__buf_4
Xfanout543 _08443_/B vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__clkbuf_8
Xfanout554 _08215_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__buf_8
Xfanout565 _07990_/B vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__buf_6
Xfanout576 _14572_/X vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__buf_8
Xfanout587 _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13199_/C1 sky130_fd_sc_hd__buf_8
X_09838_ hold3876/X _10010_/B _09837_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09838_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout598 _12513_/X vssd1 vssd1 vccd1 vccd1 _12985_/S sky130_fd_sc_hd__buf_4
XFILLER_0_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09769_ hold4761/X _10055_/B _09768_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09769_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12367_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _17090_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_213_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _17436_/D sky130_fd_sc_hd__and2_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12310_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _17067_/D sky130_fd_sc_hd__nor2_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ hold1693/X _14482_/A2 _14449_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ hold5567/X _12338_/B _11661_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11662_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ _13791_/A _13401_/B vssd1 vssd1 vccd1 vccd1 _13401_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10613_ _16695_/Q _10637_/B _10613_/C vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__and3_1
X_14381_ _15169_/A hold2413/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11593_ hold5475/X _12329_/B _11592_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16120_ _17343_/CLK _16120_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
X_10544_ hold1279/X hold3982/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13332_ _13716_/A _13332_/B vssd1 vssd1 vccd1 vccd1 _13332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16051_ _18300_/CLK _16051_/D vssd1 vssd1 vccd1 vccd1 hold708/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13263_ _13311_/A1 _13261_/X _13262_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13263_/X
+ sky130_fd_sc_hd__o211a_1
X_10475_ hold3000/X hold3882/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _15217_/A hold514/X vssd1 vssd1 vccd1 vccd1 _15002_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12214_ hold5008/X _12308_/B _12213_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _12214_/X
+ sky130_fd_sc_hd__o211a_1
X_13194_ _17575_/Q _17109_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_202_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17446_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12145_ hold3442/X _12374_/B _12144_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ hold4257/X _13871_/B _12075_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__o211a_1
X_16953_ _17860_/CLK _16953_/D vssd1 vssd1 vccd1 vccd1 _16953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_273_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18176_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15904_ _17322_/CLK _15904_/D vssd1 vssd1 vccd1 vccd1 _15904_/Q sky130_fd_sc_hd__dfxtp_1
X_11027_ hold3036/X _16833_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11028_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16884_ _18053_/CLK _16884_/D vssd1 vssd1 vccd1 vccd1 _16884_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_202_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18318_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _17726_/CLK _15835_/D vssd1 vssd1 vccd1 vccd1 _15835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _17749_/CLK _15766_/D vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12978_ _12981_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _17502_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17505_/CLK _17505_/D vssd1 vssd1 vccd1 vccd1 _17505_/Q sky130_fd_sc_hd__dfxtp_1
X_14717_ hold2172/X _14720_/B _14716_/Y _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14717_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11929_ hold5348/X _13862_/B _11928_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11929_/X
+ sky130_fd_sc_hd__o211a_1
X_15697_ _17265_/CLK _15697_/D vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17436_ _18436_/CLK _17436_/D vssd1 vssd1 vccd1 vccd1 _17436_/Q sky130_fd_sc_hd__dfxtp_1
X_14648_ _14988_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14648_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_28 _09400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_39 _14116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17370_/CLK _17367_/D vssd1 vssd1 vccd1 vccd1 _17367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14579_ hold1899/X _14610_/B _14578_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16318_ _16323_/CLK _16318_/D vssd1 vssd1 vccd1 vccd1 _16318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ _17298_/CLK _17298_/D vssd1 vssd1 vccd1 vccd1 hold803/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5007 _12208_/X vssd1 vssd1 vccd1 vccd1 _17226_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16249_ _17429_/CLK _16249_/D vssd1 vssd1 vccd1 vccd1 _16249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5018 _16967_/Q vssd1 vssd1 vccd1 vccd1 hold5018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5029 _11326_/X vssd1 vssd1 vccd1 vccd1 _16932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput102 _13121_/A vssd1 vssd1 vccd1 vccd1 hold5784/A sky130_fd_sc_hd__buf_6
XFILLER_0_179_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput113 hold5849/X vssd1 vssd1 vccd1 vccd1 hold5850/A sky130_fd_sc_hd__buf_6
Xhold4306 _12133_/X vssd1 vssd1 vccd1 vccd1 _17201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput124 hold5896/X vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_12
Xhold4317 _17141_/Q vssd1 vssd1 vccd1 vccd1 hold4317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4328 _11701_/X vssd1 vssd1 vccd1 vccd1 _17057_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput135 hold5832/X vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_12
Xoutput146 _18462_/X vssd1 vssd1 vccd1 vccd1 slv_enable sky130_fd_sc_hd__buf_12
Xhold4339 _13360_/X vssd1 vssd1 vccd1 vccd1 _17573_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3605 _11169_/Y vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3616 _10008_/Y vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3627 _17109_/Q vssd1 vssd1 vccd1 vccd1 hold3627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3638 _13854_/Y vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2904 _14085_/X vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3649 _17580_/Q vssd1 vssd1 vccd1 vccd1 hold3649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2915 _18179_/Q vssd1 vssd1 vccd1 vccd1 hold2915/X sky130_fd_sc_hd__dlygate4sd3_1
X_07953_ hold2164/X _07991_/A2 _07952_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07953_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2926 _13979_/X vssd1 vssd1 vccd1 vccd1 _17794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2937 _18038_/Q vssd1 vssd1 vccd1 vccd1 hold2937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2948 _15234_/X vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2959 _18441_/Q vssd1 vssd1 vccd1 vccd1 hold2959/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07884_ hold202/X _14789_/A vssd1 vssd1 vccd1 vccd1 _07884_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ hold3106/X _16365_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ hold1273/X _13206_/A _10580_/C vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08505_ _15509_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__or2_1
X_09485_ hold1833/X _09483_/X _09440_/X vssd1 vssd1 vccd1 vccd1 _09485_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08436_ hold2079/X _08433_/B _08435_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _08436_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_77_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18041_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _15815_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08298_ hold2300/X _08336_/A2 _08297_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _08298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5530 _11563_/X vssd1 vssd1 vccd1 vccd1 _17011_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10260_ _10998_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__or2_1
Xhold5541 _16796_/Q vssd1 vssd1 vccd1 vccd1 hold5541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5552 _10978_/X vssd1 vssd1 vccd1 vccd1 _16816_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5563 _16770_/Q vssd1 vssd1 vccd1 vccd1 hold5563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5574 _10747_/X vssd1 vssd1 vccd1 vccd1 _16739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4840 _10336_/X vssd1 vssd1 vccd1 vccd1 _16602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5585 _16782_/Q vssd1 vssd1 vccd1 vccd1 hold5585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4851 _16442_/Q vssd1 vssd1 vccd1 vccd1 hold4851/X sky130_fd_sc_hd__dlygate4sd3_1
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__or2_1
Xhold5596 _11599_/X vssd1 vssd1 vccd1 vccd1 _17023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4862 _11005_/X vssd1 vssd1 vccd1 vccd1 _16825_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4873 _16564_/Q vssd1 vssd1 vccd1 vccd1 hold4873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4884 _09958_/X vssd1 vssd1 vccd1 vccd1 _16476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4895 _16926_/Q vssd1 vssd1 vccd1 vccd1 hold4895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout340 _09369_/X vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__clkbuf_4
Xfanout351 _08721_/S vssd1 vssd1 vccd1 vccd1 _08727_/S sky130_fd_sc_hd__buf_8
XFILLER_0_233_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout362 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout373 hold513/X vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__clkbuf_8
X_13950_ hold999/X _13998_/B vssd1 vssd1 vccd1 vccd1 _13950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout384 _14734_/Y vssd1 vssd1 vccd1 vccd1 _14774_/B sky130_fd_sc_hd__buf_8
XFILLER_0_191_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout395 _14479_/B vssd1 vssd1 vccd1 vccd1 _14499_/B sky130_fd_sc_hd__buf_8
X_12901_ hold2626/X hold3161/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_199_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13881_ hold3738/X _13791_/A _13880_/X vssd1 vssd1 vccd1 vccd1 _13881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15620_ _17215_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ hold1375/X hold3355/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__or2_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12763_ hold1686/X _17432_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14502_ _15182_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14543_/B sky130_fd_sc_hd__or2_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _18272_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ hold1825/X _17062_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _11715_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15482_ _15482_/A _15482_/B vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ hold1127/X hold3760/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__mux2_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17221_/CLK _17221_/D vssd1 vssd1 vccd1 vccd1 _17221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14433_ _15547_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14433_/Y sky130_fd_sc_hd__nand2_1
X_11645_ hold1803/X hold5212/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17152_ _17280_/CLK _17152_/D vssd1 vssd1 vccd1 vccd1 _17152_/Q sky130_fd_sc_hd__dfxtp_1
Xinput15 input15/A vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_6
X_14364_ _15506_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _17979_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput26 input26/A vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_6
X_11576_ hold1650/X hold3486/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__mux2_1
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
X_16103_ _16131_/CLK _16103_/D vssd1 vssd1 vccd1 vccd1 hold685/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput48 input48/A vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_6
X_13315_ hold5268/X _12353_/B _13314_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _13315_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10527_ _10527_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17083_ _17263_/CLK _17083_/D vssd1 vssd1 vccd1 vccd1 _17083_/Q sky130_fd_sc_hd__dfxtp_1
X_14295_ hold1845/X hold756/X _14294_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _14295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ _18408_/CLK _16034_/D vssd1 vssd1 vccd1 vccd1 hold862/A sky130_fd_sc_hd__dfxtp_1
X_13246_ _13246_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13246_/X sky130_fd_sc_hd__or2_1
X_10458_ _10476_/A _10458_/B vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_454_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13177_ _13177_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__and2_1
X_10389_ _10527_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__or2_1
X_12128_ hold2538/X hold5128/X _13412_/S vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__mux2_1
X_17985_ _17985_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12059_ hold1489/X _17177_/Q _12251_/S vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__mux2_1
X_16936_ _17814_/CLK _16936_/D vssd1 vssd1 vccd1 vccd1 _16936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16867_ _18068_/CLK _16867_/D vssd1 vssd1 vccd1 vccd1 _16867_/Q sky130_fd_sc_hd__dfxtp_1
X_15818_ _17728_/CLK _15818_/D vssd1 vssd1 vccd1 vccd1 _15818_/Q sky130_fd_sc_hd__dfxtp_1
X_16798_ _17999_/CLK _16798_/D vssd1 vssd1 vccd1 vccd1 _16798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15749_ _17726_/CLK _15749_/D vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09270_ _12747_/A hold182/X vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__and2_1
XFILLER_0_111_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _15555_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08221_/X sky130_fd_sc_hd__or2_1
X_17419_ _17420_/CLK _17419_/D vssd1 vssd1 vccd1 vccd1 _17419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ _18399_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08152_ _15557_/A hold1322/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08083_ hold2424/X _08088_/B _08082_/Y _08149_/A vssd1 vssd1 vccd1 vccd1 _08083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4103 _16971_/Q vssd1 vssd1 vccd1 vccd1 hold4103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4114 _17560_/Q vssd1 vssd1 vccd1 vccd1 hold4114/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_195_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18386_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4125 _17145_/Q vssd1 vssd1 vccd1 vccd1 hold4125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4136 _13558_/X vssd1 vssd1 vccd1 vccd1 _17639_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3402 _11056_/X vssd1 vssd1 vccd1 vccd1 _16842_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4147 _17738_/Q vssd1 vssd1 vccd1 vccd1 hold4147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3413 _09607_/X vssd1 vssd1 vccd1 vccd1 _16359_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4158 _17156_/Q vssd1 vssd1 vccd1 vccd1 hold4158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4169 _16610_/Q vssd1 vssd1 vccd1 vccd1 hold4169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3424 _17593_/Q vssd1 vssd1 vccd1 vccd1 hold3424/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3435 _11977_/X vssd1 vssd1 vccd1 vccd1 _17149_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2701 _18036_/Q vssd1 vssd1 vccd1 vccd1 hold2701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3446 _17209_/Q vssd1 vssd1 vccd1 vccd1 hold3446/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3457 _11968_/X vssd1 vssd1 vccd1 vccd1 _17146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _13985_/X vssd1 vssd1 vccd1 vccd1 _17797_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08985_ hold222/X hold348/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__mux2_1
Xhold2723 _15778_/Q vssd1 vssd1 vccd1 vccd1 hold2723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3468 _17393_/Q vssd1 vssd1 vccd1 vccd1 hold3468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2734 _14462_/X vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3479 _12082_/X vssd1 vssd1 vccd1 vccd1 _17184_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2745 _16230_/Q vssd1 vssd1 vccd1 vccd1 hold2745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2756 _15106_/X vssd1 vssd1 vccd1 vccd1 _18335_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07936_ _15559_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07936_/X sky130_fd_sc_hd__or2_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2767 _15176_/X vssd1 vssd1 vccd1 vccd1 _18369_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2778 _18208_/Q vssd1 vssd1 vccd1 vccd1 hold2778/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2789 _16225_/Q vssd1 vssd1 vccd1 vccd1 hold2789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07867_ _15545_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09606_ _09984_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07798_ _07804_/A _09342_/A _09339_/B hold3163/X vssd1 vssd1 vccd1 vccd1 _07798_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_211_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ _09963_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09472_/C _09472_/D _09472_/B vssd1 vssd1 vccd1 vccd1 _09470_/C sky130_fd_sc_hd__a21o_1
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08419_ _15533_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _15559_/A _14555_/C hold329/X _09398_/X vssd1 vssd1 vccd1 vccd1 _09400_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_80_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _12204_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _11553_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6050 _16311_/Q vssd1 vssd1 vccd1 vccd1 hold6050/X sky130_fd_sc_hd__dlygate4sd3_1
X_10312_ hold3668/X _10598_/B _10311_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__o211a_1
X_13100_ hold3758/X _13099_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_105_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11292_ _12051_/A _11292_/B vssd1 vssd1 vccd1 vccd1 _11292_/X sky130_fd_sc_hd__or2_1
X_14080_ _15533_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5360 _17136_/Q vssd1 vssd1 vccd1 vccd1 hold5360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ hold922/X hold958/X _13031_/C vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__and3b_1
X_10243_ hold4803/X _10625_/B _10242_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5371 _17021_/Q vssd1 vssd1 vccd1 vccd1 hold5371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5382 _10237_/X vssd1 vssd1 vccd1 vccd1 _16569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5393 _16657_/Q vssd1 vssd1 vccd1 vccd1 hold5393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4670 _16727_/Q vssd1 vssd1 vccd1 vccd1 hold4670/X sky130_fd_sc_hd__dlygate4sd3_1
X_10174_ hold4067/X _10598_/B _10173_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _10174_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4681 _16911_/Q vssd1 vssd1 vccd1 vccd1 hold4681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4692 _12318_/Y vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3980 _16694_/Q vssd1 vssd1 vccd1 vccd1 hold3980/X sky130_fd_sc_hd__dlygate4sd3_1
X_17770_ _17834_/CLK hold248/X vssd1 vssd1 vccd1 vccd1 _17770_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3991 _10423_/X vssd1 vssd1 vccd1 vccd1 _16631_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14982_ _15523_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout170 _13808_/B vssd1 vssd1 vccd1 vccd1 _12031_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout181 _11168_/B vssd1 vssd1 vccd1 vccd1 _11738_/B sky130_fd_sc_hd__buf_4
Xfanout192 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _13886_/B sky130_fd_sc_hd__clkbuf_8
X_16721_ _18018_/CLK _16721_/D vssd1 vssd1 vccd1 vccd1 _16721_/Q sky130_fd_sc_hd__dfxtp_1
X_13933_ _13933_/A hold275/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__and2_1
XFILLER_0_135_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ _18176_/CLK _16652_/D vssd1 vssd1 vccd1 vccd1 _16652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13864_ _13864_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _17741_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_201_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _17283_/CLK _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ hold3181/X _12814_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__mux2_1
X_16583_ _18205_/CLK _16583_/D vssd1 vssd1 vccd1 vccd1 _16583_/Q sky130_fd_sc_hd__dfxtp_1
X_13795_ hold5370/X _12353_/B _13794_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _17718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18322_ _18322_/CLK hold766/X vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ hold2782/X _15547_/B _15533_/X _12657_/A vssd1 vssd1 vccd1 vccd1 _15534_/X
+ sky130_fd_sc_hd__o211a_1
X_12746_ hold3195/X _12745_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18393_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ hold665/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15465_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ hold3334/X _12676_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__mux2_1
X_17204_ _17236_/CLK _17204_/D vssd1 vssd1 vccd1 vccd1 _17204_/Q sky130_fd_sc_hd__dfxtp_1
X_14416_ hold3080/X _14446_/A2 _14415_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18184_ _18216_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _11631_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11628_/X sky130_fd_sc_hd__or2_1
X_15396_ _17343_/Q _15479_/B1 _09362_/D hold281/X vssd1 vssd1 vccd1 vccd1 _15396_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17135_ _17263_/CLK _17135_/D vssd1 vssd1 vccd1 vccd1 _17135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _15189_/A hold3232/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14348_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _11658_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold607 hold32/X vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__buf_4
Xhold618 hold618/A vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold629 hold629/A vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17066_ _17879_/CLK _17066_/D vssd1 vssd1 vccd1 vccd1 _17066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14278_ _14726_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _18422_/CLK _16017_/D vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13229_ _13228_/X hold4701/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _14567_/X vssd1 vssd1 vccd1 vccd1 _18076_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _15721_/Q vssd1 vssd1 vccd1 vccd1 hold2019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _17966_/Q vssd1 vssd1 vccd1 vccd1 hold1307/X sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ _15324_/A hold669/X vssd1 vssd1 vccd1 vccd1 _16005_/D sky130_fd_sc_hd__and2_1
Xhold1318 _18291_/Q vssd1 vssd1 vccd1 vccd1 hold1318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17968_ _17968_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1329 _16288_/Q vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16919_ _17970_/CLK _16919_/D vssd1 vssd1 vccd1 vccd1 _16919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17899_ _17899_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09322_ hold2033/X _09325_/B _09321_/Y _12969_/A vssd1 vssd1 vccd1 vccd1 _09322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ _15529_/A hold2585/X _09273_/S vssd1 vssd1 vccd1 vccd1 _09254_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ hold2791/X _08209_/B _08203_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09184_ _15513_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_376_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17696_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _08385_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__and2_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_305_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08066_ _15525_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3210 _12749_/X vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3221 _14468_/X vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3232 _17971_/Q vssd1 vssd1 vccd1 vccd1 hold3232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3243 _10002_/Y vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3254 _17508_/Q vssd1 vssd1 vccd1 vccd1 hold3254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 _16327_/Q vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2520 _18142_/Q vssd1 vssd1 vccd1 vccd1 hold2520/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2531 _16243_/Q vssd1 vssd1 vccd1 vccd1 hold2531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3276 _17509_/Q vssd1 vssd1 vccd1 vccd1 hold3276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3287 _12602_/X vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2542 _18057_/Q vssd1 vssd1 vccd1 vccd1 hold2542/X sky130_fd_sc_hd__dlygate4sd3_1
X_08968_ _15491_/A _08968_/B vssd1 vssd1 vccd1 vccd1 _16101_/D sky130_fd_sc_hd__and2_1
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3298 _12863_/X vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2553 _16172_/Q vssd1 vssd1 vccd1 vccd1 hold2553/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 _15773_/Q vssd1 vssd1 vccd1 vccd1 hold2564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 _14805_/X vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2575 _15726_/Q vssd1 vssd1 vccd1 vccd1 hold2575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1841 _18268_/Q vssd1 vssd1 vccd1 vccd1 hold1841/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ hold2399/X _07918_/B _07918_/Y _08147_/A vssd1 vssd1 vccd1 vccd1 _07919_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2586 _15590_/Q vssd1 vssd1 vccd1 vccd1 hold2586/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1852 _15212_/X vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2597 _15768_/Q vssd1 vssd1 vccd1 vccd1 hold2597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08899_ _12426_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__and2_1
Xhold1863 _18007_/Q vssd1 vssd1 vccd1 vccd1 hold1863/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_230_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1874 _13977_/X vssd1 vssd1 vccd1 vccd1 _17793_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1885 _18359_/Q vssd1 vssd1 vccd1 vccd1 hold1885/X sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ hold5020/X _11216_/B _10929_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10930_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_92_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16089_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1896 _14223_/X vssd1 vssd1 vccd1 vccd1 _17911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ hold4307/X _11147_/B _10860_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10861_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12600_ _12600_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _17376_/D sky130_fd_sc_hd__and2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13580_ hold2038/X hold3517/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ hold5517/X _11210_/B _10791_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _10792_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12531_ _12531_/A _12531_/B vssd1 vssd1 vccd1 vccd1 _17353_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _15910_/Q _15486_/A2 _09357_/B hold419/X vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _17324_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ hold2838/X _14202_/B _14200_/Y _13919_/A vssd1 vssd1 vccd1 vccd1 _14201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ hold4332/X _12365_/B _11412_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _15182_/A hold393/X vssd1 vssd1 vccd1 vccd1 _15181_/Y sky130_fd_sc_hd__nor2_2
X_12393_ hold47/X hold421/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14132_ _14758_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11344_ hold4030/X _11726_/B _11343_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11344_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14063_ hold2713/X _14107_/A2 _14062_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14063_/X
+ sky130_fd_sc_hd__o211a_1
X_11275_ hold5537/X _11753_/B _11274_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11275_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5190 _17225_/Q vssd1 vssd1 vccd1 vccd1 hold5190/X sky130_fd_sc_hd__dlygate4sd3_1
X_13014_ hold2203/X _13003_/Y _13013_/X _12531_/A vssd1 vssd1 vccd1 vccd1 _13014_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10226_ hold2170/X _16566_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__mux2_1
XTAP_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10157_ hold2246/X _16543_/Q _10613_/C vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__mux2_1
X_17822_ _17822_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ hold2006/X hold4634/X _10580_/C vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__mux2_1
X_14965_ hold2981/X _14952_/B _14964_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17753_ _17882_/CLK _17753_/D vssd1 vssd1 vccd1 vccd1 _17753_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16704_ _18228_/CLK _16704_/D vssd1 vssd1 vccd1 vccd1 _16704_/Q sky130_fd_sc_hd__dfxtp_1
X_13916_ _14758_/A hold2233/X hold124/X vssd1 vssd1 vccd1 vccd1 _13917_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_233_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17684_ _17748_/CLK _17684_/D vssd1 vssd1 vccd1 vccd1 _17684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ _14897_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14896_/Y sky130_fd_sc_hd__nor2_2
X_16635_ _18223_/CLK _16635_/D vssd1 vssd1 vccd1 vccd1 _16635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ _17736_/Q _13847_/B _13847_/C vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _18154_/CLK _16566_/D vssd1 vssd1 vccd1 vccd1 _16566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13778_ hold1910/X _17713_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18305_ _18305_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15517_ _15517_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__or2_1
X_12729_ _12738_/A _12729_/B vssd1 vssd1 vccd1 vccd1 _17419_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16497_ _18376_/CLK _16497_/D vssd1 vssd1 vccd1 vccd1 _16497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18236_ _18367_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15448_ hold546/X _15486_/A2 _15448_/B1 hold773/X vssd1 vssd1 vccd1 vccd1 _15448_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18167_ _18231_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ hold879/X _09365_/B _09392_/C hold858/X _15378_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold404 hold404/A vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ _17278_/CLK _17118_/D vssd1 vssd1 vccd1 vccd1 _17118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ _18208_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
Xhold426 hold426/A vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold437 hold437/A vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ hold5322/X _10034_/B _09939_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09940_/X
+ sky130_fd_sc_hd__o211a_1
X_17049_ _17895_/CLK _17049_/D vssd1 vssd1 vccd1 vccd1 _17049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout906 hold719/X vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__buf_8
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09871_ hold4717/X _10577_/B _09870_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09871_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 hold559/X vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__clkbuf_16
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _15213_/A vssd1 vssd1 vccd1 vccd1 _15105_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout939 _15205_/A vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__buf_12
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ hold163/X hold300/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__mux2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 la_data_in[7] vssd1 vssd1 vccd1 vccd1 hold1104/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _15722_/Q vssd1 vssd1 vccd1 vccd1 hold1115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 _15528_/X vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1137 _13924_/X vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ hold361/X _15997_/Q _08779_/S vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__mux2_1
Xhold1148 _14867_/X vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_240_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1159 _15608_/Q vssd1 vssd1 vccd1 vccd1 hold1159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _15364_/A hold483/X vssd1 vssd1 vccd1 vccd1 _15963_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09305_ hold944/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09236_ _12768_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _16229_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ hold2254/X _09164_/B _09166_/X _12909_/A vssd1 vssd1 vccd1 vccd1 _09167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08118_ _14517_/A hold1316/X hold240/X vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09098_ _15105_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ hold202/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__or2_4
XFILLER_0_222_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold971 hold979/X vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11060_ hold870/X hold3535/X _11156_/C vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__mux2_1
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3040 _09143_/X vssd1 vssd1 vccd1 vccd1 _16184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3051 _18119_/Q vssd1 vssd1 vccd1 vccd1 hold3051/X sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ _13142_/A _09933_/A _10010_/X vssd1 vssd1 vccd1 vccd1 _10011_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3062 _13965_/X vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3073 _17950_/Q vssd1 vssd1 vccd1 vccd1 hold3073/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3084 _18169_/Q vssd1 vssd1 vccd1 vccd1 hold3084/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3095 _18145_/Q vssd1 vssd1 vccd1 vccd1 hold3095/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2350 _14544_/X vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2361 _18450_/Q vssd1 vssd1 vccd1 vccd1 hold2361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2372 _14621_/X vssd1 vssd1 vccd1 vccd1 _18102_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 _08330_/X vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _09101_/X vssd1 vssd1 vccd1 vccd1 _16165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1660 _18330_/Q vssd1 vssd1 vccd1 vccd1 hold1660/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14750_ _15197_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__or2_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1671 _07882_/X vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1682 _18027_/Q vssd1 vssd1 vccd1 vccd1 hold1682/X sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ hold4579/X _12344_/B _11961_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1693 _18020_/Q vssd1 vssd1 vccd1 vccd1 hold1693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13800_/A _13701_/B vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__or2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ hold1998/X _16795_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__mux2_1
X_14681_ _14681_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14730_/B sky130_fd_sc_hd__or2_4
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ hold4445/X _13877_/B _11892_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16420_ _18363_/CLK _16420_/D vssd1 vssd1 vccd1 vccd1 _16420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13632_ _13767_/A _13632_/B vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10844_ _17973_/Q hold5477/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_298_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17858_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _18294_/CLK _16351_/D vssd1 vssd1 vccd1 vccd1 _16351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13563_ _13791_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__or2_1
X_10775_ hold3073/X _16749_/Q _11159_/C vssd1 vssd1 vccd1 vccd1 _10776_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_227_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18181_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15302_ _15489_/A _15302_/B _15302_/C _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ hold1716/X hold3250/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12514_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_180_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16282_ _18459_/CLK _16282_/D vssd1 vssd1 vccd1 vccd1 _16282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13494_ _13791_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18021_ _18052_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12445_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_212_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ hold962/X _15167_/B _15163_/Y _15032_/A vssd1 vssd1 vccd1 vccd1 hold963/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ _13888_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _17282_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14115_ hold1821/X _14142_/B _14114_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _14115_/X
+ sky130_fd_sc_hd__o211a_1
X_11327_ hold1271/X hold3831/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__mux2_1
X_15095_ _15203_/A hold734/X vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14046_ _14726_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__or2_1
X_11258_ hold3014/X hold4697/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11259_/B sky130_fd_sc_hd__mux2_1
X_10209_ _10497_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11189_ _11189_/A _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__and3_1
XFILLER_0_140_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17805_ _17808_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15997_ _18399_/CLK _15997_/D vssd1 vssd1 vccd1 vccd1 _15997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _15217_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17736_ _17736_/CLK _17736_/D vssd1 vssd1 vccd1 vccd1 _17736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14879_ hold2180/X _14882_/B _14878_/Y _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14879_/X
+ sky130_fd_sc_hd__o211a_1
X_17667_ _17667_/CLK _17667_/D vssd1 vssd1 vccd1 vccd1 _17667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _18287_/CLK _16618_/D vssd1 vssd1 vccd1 vccd1 _16618_/Q sky130_fd_sc_hd__dfxtp_1
X_17598_ _17726_/CLK _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16549_ _18233_/CLK _16549_/D vssd1 vssd1 vccd1 vccd1 _16549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09021_ _09053_/A hold573/X vssd1 vssd1 vccd1 vccd1 _16127_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18219_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5904 _09486_/X vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5915 _16313_/Q vssd1 vssd1 vccd1 vccd1 hold5915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5926 _17552_/Q vssd1 vssd1 vccd1 vccd1 hold5926/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 data_in[2] vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5937 _17546_/Q vssd1 vssd1 vccd1 vccd1 hold5937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5948 _17557_/Q vssd1 vssd1 vccd1 vccd1 hold5948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5959 data_in[16] vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 input45/X vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold256 hold35/X vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__buf_4
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold278 hold46/X vssd1 vssd1 vccd1 vccd1 input33/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_48_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_48_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_09923_ hold2250/X _16465_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__mux2_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _12396_/A vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout714 _15491_/A vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__clkbuf_4
Xfanout725 _15044_/A vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__buf_4
Xfanout736 _09063_/A vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09854_ hold1733/X _16442_/Q _10049_/C vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__mux2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout747 _08111_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout758 _13903_/A vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__buf_4
Xfanout769 fanout770/X vssd1 vssd1 vccd1 vccd1 _14538_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _13037_/A hold774/X vssd1 vssd1 vccd1 vccd1 _16021_/D sky130_fd_sc_hd__and2_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ hold1660/X hold4723/X _10601_/C vssd1 vssd1 vccd1 vccd1 _09786_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ _15454_/A hold441/X vssd1 vssd1 vccd1 vccd1 _15988_/D sky130_fd_sc_hd__and2_1
XFILLER_0_212_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ hold312/X hold413/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__mux2_1
XFILLER_0_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _12380_/A _12445_/A vssd1 vssd1 vccd1 vccd1 _08627_/S sky130_fd_sc_hd__or2_2
XFILLER_0_3_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_391_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17145_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_230_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_320_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17891_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _10560_/A _10560_/B vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ hold2347/X _09216_/B _09218_/Y _12912_/A vssd1 vssd1 vccd1 vccd1 _09219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _10533_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ hold1540/X hold4229/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12161_ hold2793/X hold5435/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11694_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12092_ hold2335/X hold4253/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__mux2_1
Xhold790 hold790/A vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _18405_/CLK _15920_/D vssd1 vssd1 vccd1 vccd1 hold907/A sky130_fd_sc_hd__dfxtp_1
X_11043_ _11139_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _17731_/CLK _15851_/D vssd1 vssd1 vccd1 vccd1 _15851_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2180 _18226_/Q vssd1 vssd1 vccd1 vccd1 hold2180/X sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ _15195_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__or2_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2191 _14323_/X vssd1 vssd1 vccd1 vccd1 _17959_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15782_ _17681_/CLK _15782_/D vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ hold2553/X _17509_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_231_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 _07941_/X vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17521_ _17523_/CLK hold923/X vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_1
X_14733_ hold2878/X _14720_/B _14732_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14733_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ hold2471/X _17139_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_408_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17886_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17481_/CLK _17452_/D vssd1 vssd1 vccd1 vccd1 _17452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _15004_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _15708_/Q hold4779/X _13862_/C vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _18346_/CLK _16403_/D vssd1 vssd1 vccd1 vccd1 _16403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13615_ hold4213/X _13814_/B _13614_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _13615_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17383_ _17459_/CLK _17383_/D vssd1 vssd1 vccd1 vccd1 _17383_/Q sky130_fd_sc_hd__dfxtp_1
X_10827_ _11667_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__or2_1
X_14595_ hold3004/X _14610_/B _14594_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16334_ _18342_/CLK _16334_/D vssd1 vssd1 vccd1 vccd1 _16334_/Q sky130_fd_sc_hd__dfxtp_1
X_13546_ hold5731/X _13832_/B _13545_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13546_/X
+ sky130_fd_sc_hd__o211a_1
X_10758_ _11052_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16265_ _17370_/CLK _16265_/D vssd1 vssd1 vccd1 vccd1 _16265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13477_ hold4569/X _13847_/B _13476_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10689_ _11553_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__or2_1
X_15216_ hold1212/X _15219_/B _15215_/Y _15024_/A vssd1 vssd1 vccd1 vccd1 _15216_/X
+ sky130_fd_sc_hd__o211a_1
X_18004_ _18064_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12428_ _12438_/A hold264/X vssd1 vssd1 vccd1 vccd1 _17307_/D sky130_fd_sc_hd__and2_1
X_16196_ _17481_/CLK _16196_/D vssd1 vssd1 vccd1 vccd1 _16196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15147_ _15201_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15147_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _17277_/Q _13868_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__and3_1
XFILLER_0_239_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3809 _09526_/X vssd1 vssd1 vccd1 vccd1 _16332_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_205_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15078_ hold1194/X _15111_/B _15077_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15078_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14029_ hold1656/X _14040_/B _14028_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _14029_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ _09954_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08521_ _08868_/B _13056_/C _17520_/Q vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_89_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17719_ _17719_/CLK _17719_/D vssd1 vssd1 vccd1 vccd1 _17719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_149_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18367_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08452_ hold999/X _08500_/B vssd1 vssd1 vccd1 vccd1 _08452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _15823_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09004_ hold215/X _16119_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5701 _17698_/Q vssd1 vssd1 vccd1 vccd1 hold5701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5712 _10096_/X vssd1 vssd1 vccd1 vccd1 _16522_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5723 _17727_/Q vssd1 vssd1 vccd1 vccd1 hold5723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5734 _13579_/X vssd1 vssd1 vccd1 vccd1 _17646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5745 _17633_/Q vssd1 vssd1 vccd1 vccd1 hold5745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5756 _13633_/X vssd1 vssd1 vccd1 vccd1 _17664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5767 hold5924/X vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5778 output87/X vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_12
Xhold5789 hold5933/X vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout500 _11093_/S vssd1 vssd1 vccd1 vccd1 _11198_/C sky130_fd_sc_hd__buf_6
XFILLER_0_228_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout511 _10400_/S vssd1 vssd1 vccd1 vccd1 _10481_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09906_ _09936_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__or2_1
Xfanout522 _09317_/B vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__buf_4
Xfanout533 _09098_/B vssd1 vssd1 vccd1 vccd1 _09118_/B sky130_fd_sc_hd__clkbuf_4
Xfanout544 _08440_/A2 vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__clkbuf_8
Xfanout555 _08173_/Y vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__buf_8
Xfanout566 _07991_/A2 vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__buf_6
X_09837_ _09933_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__or2_1
Xfanout577 hold392/X vssd1 vssd1 vccd1 vccd1 hold393/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_232_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout588 _13049_/Y vssd1 vssd1 vccd1 vccd1 _13311_/C1 sky130_fd_sc_hd__clkbuf_16
Xfanout599 _12601_/S vssd1 vssd1 vccd1 vccd1 _13000_/S sky130_fd_sc_hd__buf_6
XFILLER_0_241_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09768_ _09960_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ hold145/X hold714/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold715/A sky130_fd_sc_hd__mux2_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09963_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11730_ hold3600/X _11637_/A _11729_/X vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _12243_/A _11661_/B vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ hold2599/X hold3738/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _11194_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _16694_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_154_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14380_ _14380_/A hold659/X vssd1 vssd1 vccd1 vccd1 _17987_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11592_ _12234_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13331_ hold2083/X hold4647/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ hold5058/X _10637_/B _10542_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _10543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16050_ _16128_/CLK _16050_/D vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ _13262_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10474_ hold5126/X _10625_/B _10473_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__o211a_1
X_15001_ hold1168/X _15004_/B _15000_/Y _15070_/A vssd1 vssd1 vccd1 vccd1 _15001_/X
+ sky130_fd_sc_hd__o211a_1
X_12213_ _12213_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13193_ _13193_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__and2_1
XFILLER_0_150_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12144_ _12273_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ _12267_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__or2_1
X_16952_ _17869_/CLK _16952_/D vssd1 vssd1 vccd1 vccd1 _16952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15903_ _16126_/CLK _15903_/D vssd1 vssd1 vccd1 vccd1 hold840/A sky130_fd_sc_hd__dfxtp_1
X_11026_ hold5302/X _11216_/B _11025_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _11026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16883_ _18319_/CLK _16883_/D vssd1 vssd1 vccd1 vccd1 _16883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _17426_/CLK _15834_/D vssd1 vssd1 vccd1 vccd1 _15834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _17748_/CLK _15765_/D vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfxtp_1
X_12977_ hold3215/X _12976_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_242_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18178_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17505_/CLK _17504_/D vssd1 vssd1 vccd1 vccd1 _17504_/Q sky130_fd_sc_hd__dfxtp_1
X_14716_ _14878_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ _12024_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__or2_1
X_15696_ _17718_/CLK _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ hold3090/X _14666_/B _14646_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17435_ _17435_/CLK _17435_/D vssd1 vssd1 vccd1 vccd1 _17435_/Q sky130_fd_sc_hd__dfxtp_1
X_11859_ _12243_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _14794_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__or2_1
XANTENNA_29 _09400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _17376_/CLK _17366_/D vssd1 vssd1 vccd1 vccd1 _17366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16317_ _16320_/CLK _16317_/D vssd1 vssd1 vccd1 vccd1 _16317_/Q sky130_fd_sc_hd__dfxtp_1
X_13529_ _15815_/Q hold4934/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17297_ _17297_/CLK _17297_/D vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _17429_/CLK _16248_/D vssd1 vssd1 vccd1 vccd1 _16248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5008 _17260_/Q vssd1 vssd1 vccd1 vccd1 hold5008/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5019 _11335_/X vssd1 vssd1 vccd1 vccd1 _16935_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _13129_/A vssd1 vssd1 vccd1 vccd1 hold5782/A sky130_fd_sc_hd__buf_6
Xhold4307 _16809_/Q vssd1 vssd1 vccd1 vccd1 hold4307/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput114 hold5872/X vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_12
X_16179_ _17483_/CLK _16179_/D vssd1 vssd1 vccd1 vccd1 _16179_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput125 hold5858/X vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_12
Xhold4318 _11857_/X vssd1 vssd1 vccd1 vccd1 _17109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4329 hold6042/X vssd1 vssd1 vccd1 vccd1 hold4329/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput136 hold4585/X vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_12
Xhold3606 _17363_/Q vssd1 vssd1 vccd1 vccd1 hold3606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3617 _17561_/Q vssd1 vssd1 vccd1 vccd1 hold3617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3628 _12336_/Y vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3639 _17122_/Q vssd1 vssd1 vccd1 vccd1 hold3639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2905 _15623_/Q vssd1 vssd1 vccd1 vccd1 hold2905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2916 _14781_/X vssd1 vssd1 vccd1 vccd1 _18179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07952_ _14246_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07952_/X sky130_fd_sc_hd__or2_1
Xhold2927 _18293_/Q vssd1 vssd1 vccd1 vccd1 hold2927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2938 _14486_/X vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2949 _18163_/Q vssd1 vssd1 vccd1 vccd1 hold2949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07883_ hold689/X hold764/A hold732/X hold752/X vssd1 vssd1 vccd1 vccd1 _14789_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09622_ hold5399/X _10034_/B _09621_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09553_ hold4755/X _10055_/B _09552_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08504_ hold203/X _14897_/A vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__or2_2
XFILLER_0_194_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09484_ _09483_/X _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _16322_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_148_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08435_ _14328_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ hold1016/X _15815_/Q hold134/X vssd1 vssd1 vccd1 vccd1 _08366_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ _14246_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08297_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5520 _11296_/X vssd1 vssd1 vccd1 vccd1 _16922_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5531 _17086_/Q vssd1 vssd1 vccd1 vccd1 hold5531/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5542 _10822_/X vssd1 vssd1 vccd1 vccd1 _16764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5553 _16893_/Q vssd1 vssd1 vccd1 vccd1 hold5553/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5564 _10744_/X vssd1 vssd1 vccd1 vccd1 _16738_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4830 _10339_/X vssd1 vssd1 vccd1 vccd1 _16603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5575 _17013_/Q vssd1 vssd1 vccd1 vccd1 hold5575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4841 _16416_/Q vssd1 vssd1 vccd1 vccd1 hold4841/X sky130_fd_sc_hd__dlygate4sd3_1
X_10190_ hold3063/X _16554_/Q _10190_/S vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__mux2_1
Xhold5586 _10780_/X vssd1 vssd1 vccd1 vccd1 _16750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4852 _09760_/X vssd1 vssd1 vccd1 vccd1 _16410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5597 _16466_/Q vssd1 vssd1 vccd1 vccd1 hold5597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4863 _16699_/Q vssd1 vssd1 vccd1 vccd1 hold4863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4874 _10126_/X vssd1 vssd1 vccd1 vccd1 _16532_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4885 _16660_/Q vssd1 vssd1 vccd1 vccd1 hold4885/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout330 _10542_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__buf_4
Xhold4896 _11787_/Y vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout341 _09368_/Y vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__clkbuf_8
Xfanout352 _08685_/S vssd1 vssd1 vccd1 vccd1 _08721_/S sky130_fd_sc_hd__buf_8
XFILLER_0_195_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout363 _15171_/B vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__buf_8
XFILLER_0_233_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout374 _14958_/B vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__buf_6
Xfanout385 _14734_/Y vssd1 vssd1 vccd1 vccd1 _14772_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout396 _14487_/B vssd1 vssd1 vccd1 vccd1 _14482_/A2 sky130_fd_sc_hd__buf_6
X_12900_ _12909_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _17476_/D sky130_fd_sc_hd__and2_1
X_13880_ _17747_/Q _13880_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__and3_1
XFILLER_0_198_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _12912_/A _12831_/B vssd1 vssd1 vccd1 vccd1 _17453_/D sky130_fd_sc_hd__and2_1
XFILLER_0_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15550_ hold2134/X _15547_/B _15549_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _15550_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12768_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _17430_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ _15182_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14501_/Y sky130_fd_sc_hd__nor2_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ hold3833/X _12308_/B _11712_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__o211a_1
X_15481_ _15481_/A1 _15474_/X _15480_/X _15481_/B1 hold5892/A vssd1 vssd1 vccd1 vccd1
+ _15481_/X sky130_fd_sc_hd__a32o_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12693_ _12696_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _17407_/D sky130_fd_sc_hd__and2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ hold911/X _14433_/B _14431_/Y _14366_/A vssd1 vssd1 vccd1 vccd1 hold912/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17897_/CLK _17220_/D vssd1 vssd1 vccd1 vccd1 _17220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11644_ hold5220/X _11738_/B _11643_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11644_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17151_ _17903_/CLK _17151_/D vssd1 vssd1 vccd1 vccd1 _17151_/Q sky130_fd_sc_hd__dfxtp_1
X_14363_ _15205_/A hold1056/X hold333/X vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__mux2_1
Xinput16 input16/A vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_11575_ hold5648/X _11789_/B _11574_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__o211a_1
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
X_16102_ _18423_/CLK _16102_/D vssd1 vssd1 vccd1 vccd1 hold678/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
X_13314_ _13794_/A _13314_/B vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__or2_1
X_10526_ hold1773/X _16666_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput49 input49/A vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
X_17082_ _17862_/CLK _17082_/D vssd1 vssd1 vccd1 vccd1 _17082_/Q sky130_fd_sc_hd__dfxtp_1
X_14294_ _14974_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16033_ _18403_/CLK _16033_/D vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__dfxtp_1
X_13245_ _13244_/X hold4621/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__mux2_1
X_10457_ hold1579/X _16643_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _13169_/X _13175_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17540_/D sky130_fd_sc_hd__o21a_1
X_10388_ hold2524/X _16620_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ hold5389/X _12353_/B _12126_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17984_ _17985_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 hold645/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12058_ hold4551/X _12344_/B _12057_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _12058_/X
+ sky130_fd_sc_hd__o211a_1
X_16935_ _17814_/CLK _16935_/D vssd1 vssd1 vccd1 vccd1 _16935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_423_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ hold3132/X hold5625/X _11201_/C vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__mux2_1
X_16866_ _18035_/CLK _16866_/D vssd1 vssd1 vccd1 vccd1 _16866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15817_ _17700_/CLK _15817_/D vssd1 vssd1 vccd1 vccd1 _15817_/Q sky130_fd_sc_hd__dfxtp_1
X_16797_ _18030_/CLK _16797_/D vssd1 vssd1 vccd1 vccd1 _16797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ _17254_/CLK _15748_/D vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15679_ _17171_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08220_ hold2761/X _08213_/B _08219_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17418_ _17420_/CLK _17418_/D vssd1 vssd1 vccd1 vccd1 _17418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18398_ _18398_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _15714_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17349_ _18398_/CLK _17349_/D vssd1 vssd1 vccd1 vccd1 _17349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08082_ _14946_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4104 _11347_/X vssd1 vssd1 vccd1 vccd1 _16939_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4115 _17277_/Q vssd1 vssd1 vccd1 vccd1 hold4115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4126 _11869_/X vssd1 vssd1 vccd1 vccd1 _17113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4137 _16429_/Q vssd1 vssd1 vccd1 vccd1 hold4137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4148 _13759_/X vssd1 vssd1 vccd1 vccd1 _17706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3403 _17428_/Q vssd1 vssd1 vccd1 vccd1 hold3403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3414 _17427_/Q vssd1 vssd1 vccd1 vccd1 hold3414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4159 _11902_/X vssd1 vssd1 vccd1 vccd1 _17124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3425 _13324_/X vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3436 _17146_/Q vssd1 vssd1 vccd1 vccd1 hold3436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08984_ _12438_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _16109_/D sky130_fd_sc_hd__and2_1
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2702 _14482_/X vssd1 vssd1 vccd1 vccd1 _18036_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3447 _12061_/X vssd1 vssd1 vccd1 vccd1 _17177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3458 _17682_/Q vssd1 vssd1 vccd1 vccd1 hold3458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 _17834_/Q vssd1 vssd1 vccd1 vccd1 hold2713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 _08290_/X vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3469 _12650_/X vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2735 _17897_/Q vssd1 vssd1 vccd1 vccd1 hold2735/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2746 _18325_/Q vssd1 vssd1 vccd1 vccd1 hold2746/X sky130_fd_sc_hd__dlygate4sd3_1
X_07935_ hold1425/X _07924_/B _07934_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _07935_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2757 _16178_/Q vssd1 vssd1 vccd1 vccd1 hold2757/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_164_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18375_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2768 _16198_/Q vssd1 vssd1 vccd1 vccd1 hold2768/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2779 _14841_/X vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07866_ hold2166/X _07865_/B _07865_/Y _08119_/A vssd1 vssd1 vccd1 vccd1 _07866_/X
+ sky130_fd_sc_hd__o211a_1
X_09605_ hold1638/X hold3384/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07797_ _18457_/Q _07788_/Y _18458_/Q hold3163/X _11158_/A vssd1 vssd1 vccd1 vccd1
+ _07797_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ hold2679/X _13158_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09472_/C _09472_/D _09466_/Y vssd1 vssd1 vccd1 vccd1 _16316_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ hold2158/X _08440_/A2 _08417_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09398_ hold764/X hold732/X hold531/A vssd1 vssd1 vccd1 vccd1 _09398_/X sky130_fd_sc_hd__and3_1
XFILLER_0_163_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08349_ _08349_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__and2_1
XFILLER_0_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ hold2369/X hold3934/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_6_7_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6040 la_data_in[1] vssd1 vssd1 vccd1 vccd1 hold995/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _10563_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or2_1
Xhold6051 _16317_/Q vssd1 vssd1 vccd1 vccd1 hold6051/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _17767_/Q _16921_/Q _11594_/S vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ _17520_/Q _13034_/D hold957/A vssd1 vssd1 vccd1 vccd1 hold922/A sky130_fd_sc_hd__and3_1
Xhold5350 _16398_/Q vssd1 vssd1 vccd1 vccd1 hold5350/X sky130_fd_sc_hd__dlygate4sd3_1
X_10242_ _10533_/A _10242_/B vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__or2_1
Xhold5361 _11842_/X vssd1 vssd1 vccd1 vccd1 _17104_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5372 _11497_/X vssd1 vssd1 vccd1 vccd1 _16989_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5383 _17221_/Q vssd1 vssd1 vccd1 vccd1 hold5383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5394 _10405_/X vssd1 vssd1 vccd1 vccd1 _16625_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4660 _16721_/Q vssd1 vssd1 vccd1 vccd1 hold4660/X sky130_fd_sc_hd__dlygate4sd3_1
X_10173_ _10563_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__or2_1
Xhold4671 _11190_/Y vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4682 _11742_/Y vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4693 _16735_/Q vssd1 vssd1 vccd1 vccd1 hold4693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3970 _16395_/Q vssd1 vssd1 vccd1 vccd1 hold3970/X sky130_fd_sc_hd__dlygate4sd3_1
X_14981_ hold5997/X _15004_/B hold1036/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14981_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3981 _10516_/X vssd1 vssd1 vccd1 vccd1 _16662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout160 _13808_/B vssd1 vssd1 vccd1 vccd1 _13802_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3992 _16444_/Q vssd1 vssd1 vccd1 vccd1 hold3992/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout171 fanout246/X vssd1 vssd1 vccd1 vccd1 _13808_/B sky130_fd_sc_hd__buf_4
X_16720_ _18049_/CLK _16720_/D vssd1 vssd1 vccd1 vccd1 _16720_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout182 _11150_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__clkbuf_4
Xfanout193 _12274_/A2 vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__buf_4
X_13932_ hold367/A _17772_/Q hold124/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__mux2_1
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16651_ _18262_/CLK _16651_/D vssd1 vssd1 vccd1 vccd1 _16651_/Q sky130_fd_sc_hd__dfxtp_1
X_13863_ hold4747/X _12261_/A _13862_/X vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ _17639_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12814_ hold2748/X _17449_/Q _12826_/S vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16582_ _18170_/CLK _16582_/D vssd1 vssd1 vccd1 vccd1 _16582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13794_ _13794_/A _13794_/B vssd1 vssd1 vccd1 vccd1 _13794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18321_ _18321_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _15533_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15533_/X sky130_fd_sc_hd__or2_1
X_12745_ _16246_/Q _17426_/Q _12748_/S vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__mux2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18252_ _18356_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
X_15464_ _15482_/A _15464_/B vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__and2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ hold1292/X _17403_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _14988_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__or2_1
X_17203_ _17899_/CLK _17203_/D vssd1 vssd1 vccd1 vccd1 _17203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11627_ hold2707/X hold3998/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__mux2_1
X_18183_ _18215_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
X_15395_ hold266/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17134_ _17166_/CLK _17134_/D vssd1 vssd1 vccd1 vccd1 _17134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14346_ _14350_/A _14346_/B vssd1 vssd1 vccd1 vccd1 _17970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11558_ hold3012/X hold5338/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold608 hold608/A vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _10554_/A _10509_/B vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17065_ _17815_/CLK _17065_/D vssd1 vssd1 vccd1 vccd1 _17065_/Q sky130_fd_sc_hd__dfxtp_1
Xhold619 hold619/A vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ hold1720/X _14272_/B _14276_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14277_/X
+ sky130_fd_sc_hd__o211a_1
X_11489_ hold1809/X _16987_/Q _12317_/C vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _16095_/CLK _16016_/D vssd1 vssd1 vccd1 vccd1 hold665/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13228_ hold4881/X _13227_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13159_ _13199_/A1 _13157_/X _13158_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13159_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 becStatus[3] vssd1 vssd1 vccd1 vccd1 hold929/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _17999_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1308 _14337_/X vssd1 vssd1 vccd1 vccd1 _17966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 _15015_/X vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16918_ _17935_/CLK _16918_/D vssd1 vssd1 vccd1 vccd1 _16918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17898_ _17898_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_233_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16849_ _18050_/CLK _16849_/D vssd1 vssd1 vccd1 vccd1 _16849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09321_ _15543_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09252_ _12738_/A hold945/X vssd1 vssd1 vccd1 vccd1 hold946/A sky130_fd_sc_hd__and2_1
XFILLER_0_168_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _15537_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09183_ hold1052/X _09218_/B _09182_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _09183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08134_ _15539_/A hold2386/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ hold1132/X _08097_/A2 _08064_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08065_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3200 _12740_/X vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_345_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17747_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3211 _17422_/Q vssd1 vssd1 vccd1 vccd1 hold3211/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3222 _17951_/Q vssd1 vssd1 vccd1 vccd1 hold3222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3233 _17375_/Q vssd1 vssd1 vccd1 vccd1 hold3233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3244 _17495_/Q vssd1 vssd1 vccd1 vccd1 hold3244/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2510 _17850_/Q vssd1 vssd1 vccd1 vccd1 hold2510/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3255 _12995_/X vssd1 vssd1 vccd1 vccd1 _12996_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3266 _09990_/Y vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2521 _14705_/X vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2532 _18125_/Q vssd1 vssd1 vccd1 vccd1 hold2532/X sky130_fd_sc_hd__dlygate4sd3_1
X_08967_ hold256/X hold302/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08968_/B sky130_fd_sc_hd__mux2_1
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3277 _12998_/X vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2543 _14526_/X vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3288 _17470_/Q vssd1 vssd1 vccd1 vccd1 hold3288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3299 _17469_/Q vssd1 vssd1 vccd1 vccd1 hold3299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 _09115_/X vssd1 vssd1 vccd1 vccd1 _16172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1820 _15158_/X vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2565 _08277_/X vssd1 vssd1 vccd1 vccd1 _15773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1831 _18204_/Q vssd1 vssd1 vccd1 vccd1 hold1831/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _14946_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07918_/Y sky130_fd_sc_hd__nand2_1
Xhold2576 _08180_/X vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1842 _14969_/X vssd1 vssd1 vccd1 vccd1 _18268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08898_ hold118/X hold804/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__mux2_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2587 _07893_/X vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 _18396_/Q vssd1 vssd1 vccd1 vccd1 hold1853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2598 _08267_/X vssd1 vssd1 vccd1 vccd1 _15768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1864 _14422_/X vssd1 vssd1 vccd1 vccd1 _18007_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1875 _18235_/Q vssd1 vssd1 vccd1 vccd1 hold1875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1886 _15156_/X vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07849_ _14862_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1897 _16279_/Q vssd1 vssd1 vccd1 vccd1 hold1897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ _11052_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09519_ _09987_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__or2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11658_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10791_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ hold3157/X _12529_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12530_/X sky130_fd_sc_hd__mux2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12461_ hold596/X _08597_/Y _08868_/X _12460_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold72/A sky130_fd_sc_hd__o311a_1
XFILLER_0_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ _15545_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_201_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11412_ _12246_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__or2_1
X_15180_ hold2997/X _15167_/B _15179_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _15180_/X
+ sky130_fd_sc_hd__o211a_1
X_12392_ _12436_/A _12392_/B vssd1 vssd1 vccd1 vccd1 _17289_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14131_ hold1729/X _14142_/B _14130_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _14131_/X
+ sky130_fd_sc_hd__o211a_1
X_11343_ _11631_/A _11343_/B vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14062_ _14116_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11274_ _11658_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11274_/X sky130_fd_sc_hd__or2_1
X_13013_ _15517_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__or2_1
Xhold5180 _16846_/Q vssd1 vssd1 vccd1 vccd1 hold5180/X sky130_fd_sc_hd__dlygate4sd3_1
X_10225_ hold4930/X _10631_/B _10224_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10225_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5191 _12109_/X vssd1 vssd1 vccd1 vccd1 _17193_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4490 _11053_/X vssd1 vssd1 vccd1 vccd1 _16841_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17821_ _17821_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ hold4789/X _11095_/A2 _10155_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10156_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_4
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17752_ _18405_/CLK _17752_/D vssd1 vssd1 vccd1 vccd1 _17752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10087_ hold4773/X _10571_/B _10086_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _10087_/X
+ sky130_fd_sc_hd__o211a_1
X_14964_ _15233_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ _18227_/CLK _16703_/D vssd1 vssd1 vccd1 vccd1 _16703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13915_ _13919_/A _13915_/B vssd1 vssd1 vccd1 vccd1 _17763_/D sky130_fd_sc_hd__and2_1
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17683_ _17683_/CLK _17683_/D vssd1 vssd1 vccd1 vccd1 _17683_/Q sky130_fd_sc_hd__dfxtp_1
X_14895_ hold1923/X _14882_/B _14894_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14895_/X
+ sky130_fd_sc_hd__o211a_1
X_16634_ _18222_/CLK _16634_/D vssd1 vssd1 vccd1 vccd1 _16634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13846_ _13888_/A _13846_/B vssd1 vssd1 vccd1 vccd1 _17735_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16565_ _18193_/CLK _16565_/D vssd1 vssd1 vccd1 vccd1 _16565_/Q sky130_fd_sc_hd__dfxtp_1
X_13777_ hold4507/X _13777_/A2 _13776_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10989_ _11082_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10989_/X sky130_fd_sc_hd__or2_1
X_18304_ _18373_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15516_ hold2061/X _15507_/Y _15515_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _15516_/X
+ sky130_fd_sc_hd__o211a_1
X_12728_ hold3508/X _12727_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16496_ _18389_/CLK _16496_/D vssd1 vssd1 vccd1 vccd1 _16496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18235_ _18371_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15447_ hold355/X _09392_/B _09392_/C hold304/X vssd1 vssd1 vccd1 vccd1 _15447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12659_ hold3466/X _12658_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18166_ _18166_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ hold872/X _09386_/A _15451_/A2 hold803/X vssd1 vssd1 vccd1 vccd1 _15378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17117_ _17744_/CLK _17117_/D vssd1 vssd1 vccd1 vccd1 _17117_/Q sky130_fd_sc_hd__dfxtp_1
Xhold405 hold405/A vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14329_ hold2092/X _14326_/B _14328_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14329_/X
+ sky130_fd_sc_hd__o211a_1
X_18097_ _18181_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
Xhold416 hold416/A vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold438 hold438/A vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_38_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_38_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_17048_ _17894_/CLK _17048_/D vssd1 vssd1 vccd1 vccd1 _17048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09870_ _10482_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__or2_1
Xfanout907 hold719/X vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__buf_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout918 hold559/X vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_239_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 hold1084/X vssd1 vssd1 vccd1 vccd1 hold1085/A sky130_fd_sc_hd__buf_6
X_08821_ _12416_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _16029_/D sky130_fd_sc_hd__and2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1105 hold1105/A vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _08168_/X vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _15344_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _15996_/D sky130_fd_sc_hd__and2_1
Xhold1127 _16229_/Q vssd1 vssd1 vccd1 vccd1 hold1127/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1138 _15859_/Q vssd1 vssd1 vccd1 vccd1 hold1138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 la_data_in[0] vssd1 vssd1 vccd1 vccd1 hold1149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ hold163/X hold482/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold483/A sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ hold3100/X _09325_/B _09303_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ hold999/X hold1127/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09166_ _15549_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ _08117_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09097_ hold3065/X _09106_/B _09096_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08048_ hold202/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08048_/Y sky130_fd_sc_hd__nor2_2
Xhold950 hold950/A vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_222_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__clkbuf_16
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3030 _15140_/X vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10010_ _16494_/Q _10010_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__and3_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3041 _18006_/Q vssd1 vssd1 vccd1 vccd1 hold3041/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3052 _14657_/X vssd1 vssd1 vccd1 vccd1 _18119_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3063 _18110_/Q vssd1 vssd1 vccd1 vccd1 hold3063/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _13110_/A _09987_/A _09998_/X vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__a21oi_1
Xhold3074 _14305_/X vssd1 vssd1 vccd1 vccd1 _17950_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 _14729_/X vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3085 _14761_/X vssd1 vssd1 vccd1 vccd1 _18169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3096 _14711_/X vssd1 vssd1 vccd1 vccd1 _18145_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 _17932_/Q vssd1 vssd1 vccd1 vccd1 hold2351/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2362 _15548_/X vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 _15785_/Q vssd1 vssd1 vccd1 vccd1 hold2373/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2384 _15688_/Q vssd1 vssd1 vccd1 vccd1 hold2384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1650 _17862_/Q vssd1 vssd1 vccd1 vccd1 hold1650/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 _16192_/Q vssd1 vssd1 vccd1 vccd1 hold2395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1661 _15096_/X vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _12057_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__or2_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1672 _18249_/Q vssd1 vssd1 vccd1 vccd1 hold1672/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1683 _14464_/X vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 _14450_/X vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ hold5611/X _11768_/B _10911_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _10912_/X
+ sky130_fd_sc_hd__o211a_1
X_13700_ hold2597/X _17687_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13701_/B sky130_fd_sc_hd__mux2_1
X_14680_ _14681_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14680_/Y sky130_fd_sc_hd__nor2_2
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11892_ _13782_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13631_ hold1395/X hold5747/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10843_ hold5607/X _11216_/B _10842_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10843_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _18293_/CLK _16350_/D vssd1 vssd1 vccd1 vccd1 _16350_/Q sky130_fd_sc_hd__dfxtp_1
X_13562_ hold1260/X hold4243/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10774_ hold5336/X _11159_/B _10773_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _10774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15301_ _16294_/Q _15477_/A2 _15487_/B1 hold832/X _15300_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/D sky130_fd_sc_hd__a221o_1
X_12513_ _13048_/A hold2124/X _07809_/X _07789_/A vssd1 vssd1 vccd1 vccd1 _12513_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16281_ _18460_/CLK _16281_/D vssd1 vssd1 vccd1 vccd1 _16281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ hold1128/X _17618_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18020_ _18052_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
X_15232_ hold1853/X _15219_/B _15231_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__o211a_1
X_12444_ _12444_/A hold416/X vssd1 vssd1 vccd1 vccd1 _17315_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_267_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18026_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15163_ _15217_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__nand2_1
X_12375_ hold3639/X _13461_/A _12374_/X vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14114_ _14794_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11326_ hold5028/X _11617_/A2 _11325_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__o211a_1
X_15094_ hold3193/X _15113_/B _15093_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15094_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ hold1549/X _14038_/B _14044_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ hold5411/X _11732_/B _11256_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _11257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10208_ hold2498/X _16560_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11188_ _11218_/A _11188_/B vssd1 vssd1 vccd1 vccd1 _16886_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ _17804_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10139_ hold2405/X hold4701/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__mux2_1
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _18408_/CLK _15996_/D vssd1 vssd1 vccd1 vccd1 hold866/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17735_ _17745_/CLK _17735_/D vssd1 vssd1 vccd1 vccd1 _17735_/Q sky130_fd_sc_hd__dfxtp_1
X_14947_ hold2490/X _14946_/B _14946_/Y _15158_/C1 vssd1 vssd1 vccd1 vccd1 _14947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17666_ _17666_/CLK _17666_/D vssd1 vssd1 vccd1 vccd1 _17666_/Q sky130_fd_sc_hd__dfxtp_1
X_14878_ _14878_/A _14882_/B vssd1 vssd1 vccd1 vccd1 _14878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_216_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _18201_/CLK _16617_/D vssd1 vssd1 vccd1 vccd1 _16617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13829_ _17730_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__and3_1
XFILLER_0_147_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17597_ _17722_/CLK _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16548_ _18234_/CLK _16548_/D vssd1 vssd1 vccd1 vccd1 _16548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _18294_/CLK _16479_/D vssd1 vssd1 vccd1 vccd1 _16479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09020_ hold98/X _16127_/Q _09062_/S vssd1 vssd1 vccd1 vccd1 hold573/A sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18218_ _18230_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5905 _16175_/Q vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__buf_1
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18149_ _18181_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5916 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold5916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__buf_4
Xhold5927 _17551_/Q vssd1 vssd1 vccd1 vccd1 hold5927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5938 _17545_/Q vssd1 vssd1 vccd1 vccd1 hold5938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold94/X vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5949 _17529_/Q vssd1 vssd1 vccd1 vccd1 hold5949/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__buf_4
XFILLER_0_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 input33/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09922_ hold5198/X _10034_/B _09921_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09922_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout704 _12396_/A vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__buf_4
XFILLER_0_106_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout715 _15491_/A vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout726 _15044_/A vssd1 vssd1 vccd1 vccd1 _15032_/A sky130_fd_sc_hd__buf_4
X_09853_ hold3345/X _10007_/B _09852_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09853_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout737 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__buf_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _08111_/A vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__buf_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _13903_/A vssd1 vssd1 vccd1 vccd1 _08117_/A sky130_fd_sc_hd__buf_4
XFILLER_0_226_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ hold554/X hold773/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold774/A sky130_fd_sc_hd__mux2_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ hold5032/X _10070_/B _09783_/X _09976_/C1 vssd1 vssd1 vccd1 vccd1 _09784_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ hold215/X hold440/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold441/A sky130_fd_sc_hd__mux2_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _12531_/A hold642/X vssd1 vssd1 vccd1 vccd1 _15954_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08597_ _17519_/Q _17518_/Q vssd1 vssd1 vccd1 vccd1 _08597_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09218_ _15547_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10490_ hold1801/X hold5240/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_360_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17178_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09149_ hold2221/X _09164_/B _09148_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09149_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ hold4110/X _13868_/B _12159_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _12160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11111_ hold2323/X hold4467/X _11768_/C vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12091_ hold3480/X _13877_/B _12090_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _12091_/X
+ sky130_fd_sc_hd__o211a_1
Xhold780 hold780/A vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 hold791/A vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ hold2620/X hold3444/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__mux2_1
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _17613_/CLK _15850_/D vssd1 vssd1 vccd1 vccd1 _15850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2170 _18122_/Q vssd1 vssd1 vccd1 vccd1 hold2170/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2181 _14879_/X vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14801_ hold2862/X _14828_/B _14800_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14801_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _15643_/Q vssd1 vssd1 vccd1 vccd1 hold2192/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _17739_/CLK _15781_/D vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12996_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _17507_/D sky130_fd_sc_hd__and2_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17520_ _17523_/CLK _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1480 _14975_/X vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1491 _18257_/Q vssd1 vssd1 vccd1 vccd1 hold1491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _15233_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__or2_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ hold4160/X _12347_/B _11943_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17481_/CLK _17451_/D vssd1 vssd1 vccd1 vccd1 _17451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ hold2170/X _14666_/B _14662_/Y _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14663_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11875_ hold5461/X _12353_/B _11874_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _18351_/CLK _16402_/D vssd1 vssd1 vccd1 vccd1 _16402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _13800_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13614_/X sky130_fd_sc_hd__or2_1
X_10826_ hold2899/X _16766_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _10827_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17382_ _17459_/CLK _17382_/D vssd1 vssd1 vccd1 vccd1 _17382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ _14988_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14594_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_448_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17189_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ _18276_/CLK _16333_/D vssd1 vssd1 vccd1 vccd1 _16333_/Q sky130_fd_sc_hd__dfxtp_1
X_10757_ hold1883/X _16743_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__mux2_1
X_13545_ _13767_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _17376_/CLK _16264_/D vssd1 vssd1 vccd1 vccd1 _16264_/Q sky130_fd_sc_hd__dfxtp_1
X_13476_ _13746_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10688_ hold2636/X hold3604/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _18003_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
X_12427_ hold263/X _17307_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__mux2_1
X_15215_ _15215_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16195_ _17481_/CLK _16195_/D vssd1 vssd1 vccd1 vccd1 _16195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15146_ hold1996/X _15165_/B _15145_/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 _15146_/X
+ sky130_fd_sc_hd__o211a_1
X_12358_ _13825_/A _12358_/B vssd1 vssd1 vccd1 vccd1 _17276_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11309_ hold2060/X _16927_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__mux2_1
X_15077_ _15131_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12289_ hold3845/X _12293_/B _12288_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12289_/X
+ sky130_fd_sc_hd__o211a_1
X_14028_ _15535_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15979_ _17298_/CLK _15979_/D vssd1 vssd1 vccd1 vccd1 hold879/A sky130_fd_sc_hd__dfxtp_1
X_08520_ _18458_/Q _13057_/B vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_222_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17718_ _17718_/CLK _17718_/D vssd1 vssd1 vccd1 vccd1 _17718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08451_ hold1312/X _08488_/B _08450_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _15854_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17649_ _17681_/CLK _17649_/D vssd1 vssd1 vccd1 vccd1 _17649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _14330_/A hold1006/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_189_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17525_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ _09053_/A hold373/X vssd1 vssd1 vccd1 vccd1 _16118_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5702 _13639_/X vssd1 vssd1 vccd1 vccd1 _17666_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5713 _17695_/Q vssd1 vssd1 vccd1 vccd1 hold5713/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5724 _13726_/X vssd1 vssd1 vccd1 vccd1 _17695_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5735 _17603_/Q vssd1 vssd1 vccd1 vccd1 hold5735/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5746 _13444_/X vssd1 vssd1 vccd1 vccd1 _17601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5757 _17614_/Q vssd1 vssd1 vccd1 vccd1 hold5757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5768 output79/X vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_83_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5779 hold5929/X vssd1 vssd1 vccd1 vccd1 _13137_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout501 _11093_/S vssd1 vssd1 vccd1 vccd1 _11216_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ hold1835/X _16459_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__mux2_1
Xfanout512 _10589_/C vssd1 vssd1 vccd1 vccd1 _10625_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout523 _09338_/A2 vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__buf_4
Xfanout534 _09066_/Y vssd1 vssd1 vccd1 vccd1 _09119_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout545 _08393_/Y vssd1 vssd1 vccd1 vccd1 _08440_/A2 sky130_fd_sc_hd__buf_8
Xfanout556 _08173_/Y vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__buf_6
X_09836_ hold1076/X _16436_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__mux2_1
Xfanout567 _07938_/Y vssd1 vssd1 vccd1 vccd1 _07991_/A2 sky130_fd_sc_hd__buf_8
Xfanout578 _14163_/B vssd1 vssd1 vccd1 vccd1 _14502_/B sky130_fd_sc_hd__buf_6
Xfanout589 _12751_/S vssd1 vssd1 vccd1 vccd1 _12763_/S sky130_fd_sc_hd__buf_6
XFILLER_0_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ hold2208/X _16413_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _12412_/A hold817/X vssd1 vssd1 vccd1 vccd1 _15980_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ hold1460/X hold4020/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__mux2_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ hold222/X hold643/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold644/A sky130_fd_sc_hd__mux2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ hold1468/X hold5545/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__mux2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10611_ hold3581/X _10497_/A _10610_/X vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11591_ hold1729/X hold5371/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13330_ hold3417/X _13802_/B _13329_/X _13714_/C1 vssd1 vssd1 vccd1 vccd1 _13330_/X
+ sky130_fd_sc_hd__o211a_1
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13261_ _13260_/X hold4639/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10473_ _10533_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ _15215_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12212_ hold1746/X _17228_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__mux2_1
X_13192_ _13185_/X _13191_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17542_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12143_ hold1373/X _17205_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12074_ hold1563/X hold4071/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__mux2_1
X_16951_ _17902_/CLK _16951_/D vssd1 vssd1 vccd1 vccd1 _16951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15902_ _16097_/CLK _15902_/D vssd1 vssd1 vccd1 vccd1 hold342/A sky130_fd_sc_hd__dfxtp_1
X_11025_ _11121_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _18019_/CLK _16882_/D vssd1 vssd1 vccd1 vccd1 _16882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _17723_/CLK _15833_/D vssd1 vssd1 vccd1 vccd1 _15833_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _17683_/CLK _15764_/D vssd1 vssd1 vccd1 vccd1 _15764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ hold2025/X _17503_/Q _12985_/S vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17879_/CLK _17503_/D vssd1 vssd1 vccd1 vccd1 _17503_/Q sky130_fd_sc_hd__dfxtp_1
X_14715_ hold1642/X _14714_/B _14714_/Y _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14715_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11927_ hold2592/X _17133_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15695_ _17769_/CLK _15695_/D vssd1 vssd1 vccd1 vccd1 _15695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17434_ _17435_/CLK _17434_/D vssd1 vssd1 vccd1 vccd1 _17434_/Q sky130_fd_sc_hd__dfxtp_1
X_14646_ _15201_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__or2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ hold2552/X hold4952/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_282_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17365_ _17365_/CLK _17365_/D vssd1 vssd1 vccd1 vccd1 _17365_/Q sky130_fd_sc_hd__dfxtp_1
X_10809_ _11100_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
XANTENNA_19 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14577_ hold1346/X _14612_/B _14576_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11789_ _17087_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_211_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18362_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16316_ _16323_/CLK _16316_/D vssd1 vssd1 vccd1 vccd1 _16316_/Q sky130_fd_sc_hd__dfxtp_1
X_13528_ hold3866/X _13814_/B _13527_/X _13720_/C1 vssd1 vssd1 vccd1 vccd1 _13528_/X
+ sky130_fd_sc_hd__o211a_1
X_17296_ _18402_/CLK _17296_/D vssd1 vssd1 vccd1 vccd1 hold574/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16247_ _17425_/CLK _16247_/D vssd1 vssd1 vccd1 vccd1 _16247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13459_ hold4348/X _13847_/B _13458_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5009 _12214_/X vssd1 vssd1 vccd1 vccd1 _17228_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput104 _18461_/X vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_12
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4308 _10861_/X vssd1 vssd1 vccd1 vccd1 _16777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput115 hold5894/X vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_12
X_16178_ _17483_/CLK _16178_/D vssd1 vssd1 vccd1 vccd1 _16178_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4319 _17025_/Q vssd1 vssd1 vccd1 vccd1 hold4319/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput126 hold5864/X vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_12
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput137 hold5846/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_12
X_15129_ _15183_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3607 _16546_/Q vssd1 vssd1 vccd1 vccd1 hold3607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3618 _13803_/Y vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3629 _17583_/Q vssd1 vssd1 vccd1 vccd1 hold3629/X sky130_fd_sc_hd__dlygate4sd3_1
X_07951_ hold1563/X _07991_/A2 _07950_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07951_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2906 _07961_/X vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2917 _18032_/Q vssd1 vssd1 vccd1 vccd1 hold2917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2928 _15019_/X vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2939 _17817_/Q vssd1 vssd1 vccd1 vccd1 hold2939/X sky130_fd_sc_hd__dlygate4sd3_1
X_07882_ hold1670/X _07865_/B _07881_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _07882_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09621_ _09843_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ _09960_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09552_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ hold203/X _14897_/A vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nor2_2
X_09483_ hold895/X hold850/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and3_1
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ hold2588/X _08433_/B _08433_/Y _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ _12750_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _15814_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ hold1192/X _08336_/A2 _08295_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5510 _11272_/X vssd1 vssd1 vccd1 vccd1 _16914_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5521 _16850_/Q vssd1 vssd1 vccd1 vccd1 hold5521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5532 _11692_/X vssd1 vssd1 vccd1 vccd1 _17054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5543 _16837_/Q vssd1 vssd1 vccd1 vccd1 hold5543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5554 _11113_/X vssd1 vssd1 vccd1 vccd1 _16861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4820 _09658_/X vssd1 vssd1 vccd1 vccd1 _16376_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5565 _16892_/Q vssd1 vssd1 vccd1 vccd1 hold5565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4831 _16503_/Q vssd1 vssd1 vccd1 vccd1 hold4831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5576 _11473_/X vssd1 vssd1 vccd1 vccd1 _16981_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4842 _09682_/X vssd1 vssd1 vccd1 vccd1 _16384_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5587 _16984_/Q vssd1 vssd1 vccd1 vccd1 hold5587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4853 _16668_/Q vssd1 vssd1 vccd1 vccd1 hold4853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17517_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5598 _09832_/X vssd1 vssd1 vccd1 vccd1 _16434_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4864 _10531_/X vssd1 vssd1 vccd1 vccd1 _16667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4875 _16651_/Q vssd1 vssd1 vccd1 vccd1 hold4875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4886 _10414_/X vssd1 vssd1 vccd1 vccd1 _16628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout320 fanout334/X vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4897 _16581_/Q vssd1 vssd1 vccd1 vccd1 hold4897/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_6_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17878_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout331 _10542_/A vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__buf_4
Xfanout342 _09368_/Y vssd1 vssd1 vccd1 vccd1 _15480_/A sky130_fd_sc_hd__buf_4
Xfanout353 _08655_/S vssd1 vssd1 vccd1 vccd1 _08661_/S sky130_fd_sc_hd__buf_8
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout364 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15167_/B sky130_fd_sc_hd__buf_8
Xfanout375 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__buf_8
Xfanout386 _14730_/B vssd1 vssd1 vccd1 vccd1 _14732_/B sky130_fd_sc_hd__buf_6
XFILLER_0_198_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09819_ _09933_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__or2_1
Xfanout397 _14447_/Y vssd1 vssd1 vccd1 vccd1 _14487_/B sky130_fd_sc_hd__buf_8
XFILLER_0_92_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ hold3353/X _12829_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_201_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12761_ hold3730/X _12760_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__mux2_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ hold870/X _14487_/B _14499_/X _14368_/A vssd1 vssd1 vccd1 vccd1 hold871/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11712_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__or2_1
X_15480_ _15480_/A _15480_/B _15480_/C _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_167_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12692_ hold4242/X _12691_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14431_ _15219_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__nand2_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11643_ _11643_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17150_ _17278_/CLK _17150_/D vssd1 vssd1 vccd1 vccd1 _17150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14362_ _14362_/A _14362_/B vssd1 vssd1 vccd1 vccd1 _17978_/D sky130_fd_sc_hd__and2_1
X_11574_ _11670_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 input17/A vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_6
XFILLER_0_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_6
X_16101_ _18411_/CLK _16101_/D vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10525_ hold5140/X _10619_/B _10524_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10525_/X
+ sky130_fd_sc_hd__o211a_1
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
X_13313_ hold1320/X _17558_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14293_ hold1883/X hold756/X _14292_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _14293_/X
+ sky130_fd_sc_hd__o211a_1
X_17081_ _17767_/CLK _17081_/D vssd1 vssd1 vccd1 vccd1 _17081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16032_ _16077_/CLK _16032_/D vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__dfxtp_1
X_13244_ hold4960/X _13243_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__mux2_2
X_10456_ hold3916/X _10646_/B _10455_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13175_ _13199_/A1 _13173_/X _13174_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13175_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_62_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10387_ hold4875/X _10577_/B _10386_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12126_ _13794_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17983_ _18016_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
X_12057_ _12057_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__or2_1
X_16934_ _17875_/CLK _16934_/D vssd1 vssd1 vccd1 vccd1 _16934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ hold5318/X _11198_/B _11007_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16865_ _17970_/CLK _16865_/D vssd1 vssd1 vccd1 vccd1 _16865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15816_ _17730_/CLK _15816_/D vssd1 vssd1 vccd1 vccd1 _15816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16796_ _17997_/CLK _16796_/D vssd1 vssd1 vccd1 vccd1 _16796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_463_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17431_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15747_ _17590_/CLK _15747_/D vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ hold3283/X _12958_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12959_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15678_ _17170_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17417_ _17420_/CLK _17417_/D vssd1 vssd1 vccd1 vccd1 _17417_/Q sky130_fd_sc_hd__dfxtp_1
X_14629_ hold1813/X _14664_/B _14628_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14629_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18397_ _18397_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _14782_/A hold2117/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17348_ _17517_/CLK _17348_/D vssd1 vssd1 vccd1 vccd1 _17348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08081_ hold2428/X _08088_/B _08080_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _17903_/CLK _17279_/D vssd1 vssd1 vccd1 vccd1 _17279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4105 _16767_/Q vssd1 vssd1 vccd1 vccd1 hold4105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4116 _12265_/X vssd1 vssd1 vccd1 vccd1 _17245_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4127 _17268_/Q vssd1 vssd1 vccd1 vccd1 hold4127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4138 _09721_/X vssd1 vssd1 vccd1 vccd1 _16397_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3404 _12755_/X vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4149 _17689_/Q vssd1 vssd1 vccd1 vccd1 hold4149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3415 _17382_/Q vssd1 vssd1 vccd1 vccd1 hold3415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3426 _16365_/Q vssd1 vssd1 vccd1 vccd1 hold3426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3437 _11872_/X vssd1 vssd1 vccd1 vccd1 _17114_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08983_ hold578/X hold592/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__mux2_1
Xhold2703 _18084_/Q vssd1 vssd1 vccd1 vccd1 hold2703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3448 _17273_/Q vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2714 _14063_/X vssd1 vssd1 vccd1 vccd1 _17834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3459 _13591_/X vssd1 vssd1 vccd1 vccd1 _17650_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 _17846_/Q vssd1 vssd1 vccd1 vccd1 hold2725/X sky130_fd_sc_hd__dlygate4sd3_1
X_07934_ _15557_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__or2_1
Xhold2736 _14193_/X vssd1 vssd1 vccd1 vccd1 _17897_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2747 _15086_/X vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _09131_/X vssd1 vssd1 vccd1 vccd1 _16178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 _09171_/X vssd1 vssd1 vccd1 vccd1 _16198_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _14878_/A _07865_/B vssd1 vssd1 vccd1 vccd1 _07865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_223_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09604_ hold4020/X _10004_/B _09603_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09604_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07796_ _11158_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_196_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09535_ hold3843/X _10019_/B _09534_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09535_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_133_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17347_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09472_/C _09472_/D _09484_/B vssd1 vssd1 vccd1 vccd1 _09466_/Y sky130_fd_sc_hd__o21ai_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _15531_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__or2_1
X_09397_ hold5866/A _09342_/B _09342_/Y _09396_/X _12404_/A vssd1 vssd1 vccd1 vccd1
+ _09397_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _14403_/A hold2053/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08279_ hold1622/X _08268_/B _08278_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6030 la_data_in[5] vssd1 vssd1 vccd1 vccd1 hold522/A sky130_fd_sc_hd__dlygate4sd3_1
X_10310_ hold2492/X _16594_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__mux2_1
Xhold6041 _16313_/Q vssd1 vssd1 vccd1 vccd1 hold6041/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6052 data_in[14] vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ hold5569/X _11768_/B _11289_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5340 _17264_/Q vssd1 vssd1 vccd1 vccd1 hold5340/X sky130_fd_sc_hd__dlygate4sd3_1
X_10241_ hold2774/X hold3677/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__mux2_1
Xhold5351 _09628_/X vssd1 vssd1 vccd1 vccd1 _16366_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5362 _16426_/Q vssd1 vssd1 vccd1 vccd1 hold5362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5373 _16622_/Q vssd1 vssd1 vccd1 vccd1 hold5373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5384 _12097_/X vssd1 vssd1 vccd1 vccd1 _17189_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4650 _10638_/Y vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5395 _16940_/Q vssd1 vssd1 vccd1 vccd1 hold5395/X sky130_fd_sc_hd__dlygate4sd3_1
X_10172_ hold3047/X _16548_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__mux2_1
Xhold4661 _11172_/Y vssd1 vssd1 vccd1 vccd1 _11173_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4672 _17097_/Q vssd1 vssd1 vccd1 vccd1 hold4672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4683 _16903_/Q vssd1 vssd1 vccd1 vccd1 hold4683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4694 _11214_/Y vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3960 _16366_/Q vssd1 vssd1 vccd1 vccd1 hold3960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3971 _09619_/X vssd1 vssd1 vccd1 vccd1 _16363_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14980_ _15195_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_233_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3982 _16672_/Q vssd1 vssd1 vccd1 vccd1 hold3982/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout150 _12974_/S vssd1 vssd1 vccd1 vccd1 _12749_/S sky130_fd_sc_hd__buf_4
Xhold3993 _09766_/X vssd1 vssd1 vccd1 vccd1 _16412_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout161 _13808_/B vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__buf_4
Xfanout172 _11617_/A2 vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__buf_4
XFILLER_0_195_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout183 fanout246/X vssd1 vssd1 vccd1 vccd1 _11150_/B sky130_fd_sc_hd__buf_4
X_13931_ _13933_/A hold125/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__and2_1
Xfanout194 _12274_/A2 vssd1 vssd1 vccd1 vccd1 _13877_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16650_ _18052_/CLK _16650_/D vssd1 vssd1 vccd1 vccd1 _16650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13862_ _17741_/Q _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15601_ _17237_/CLK _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _12912_/A _12813_/B vssd1 vssd1 vccd1 vccd1 _17447_/D sky130_fd_sc_hd__and2_1
XFILLER_0_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16581_ _18201_/CLK _16581_/D vssd1 vssd1 vccd1 vccd1 _16581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13793_ hold2772/X hold5238/X _13793_/S vssd1 vssd1 vccd1 vccd1 _13794_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18320_ _18384_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ hold2566/X _15547_/B _15531_/X _12654_/A vssd1 vssd1 vccd1 vccd1 _15532_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12750_/A _12744_/B vssd1 vssd1 vccd1 vccd1 _17424_/D sky130_fd_sc_hd__and2_1
XFILLER_0_195_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18321_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15481_/A1 _15455_/X _15462_/X _15481_/B1 _18420_/Q vssd1 vssd1 vccd1 vccd1
+ _15463_/X sky130_fd_sc_hd__a32o_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12810_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _17401_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17202_ _17266_/CLK _17202_/D vssd1 vssd1 vccd1 vccd1 _17202_/Q sky130_fd_sc_hd__dfxtp_1
X_14414_ hold3124/X _14446_/A2 _14413_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _14414_/X
+ sky130_fd_sc_hd__o211a_1
X_18182_ _18182_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ hold5224/X _12299_/B _11625_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11626_/X
+ sky130_fd_sc_hd__o211a_1
X_15394_ _15394_/A _15394_/B vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_231_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17133_ _17198_/CLK _17133_/D vssd1 vssd1 vccd1 vccd1 _17133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14345_ _14794_/A hold1741/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14346_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ hold5294/X _12314_/B _11556_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10508_ hold1791/X _16660_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10509_/B sky130_fd_sc_hd__mux2_1
Xhold609 hold609/A vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _17129_/CLK _17064_/D vssd1 vssd1 vccd1 vccd1 _17064_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_28_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_28_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14276_ _14330_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or2_1
X_11488_ hold5501/X _12338_/B _11487_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _11488_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16015_ _18422_/CLK _16015_/D vssd1 vssd1 vccd1 vccd1 _16015_/Q sky130_fd_sc_hd__dfxtp_1
X_10439_ hold3025/X hold5000/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__mux2_1
X_13227_ _13226_/X _16921_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13227_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13158_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__or2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ hold5190/X _12299_/B _12108_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _12109_/X
+ sky130_fd_sc_hd__o211a_1
X_13089_ _13089_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__and2_1
X_17966_ _17966_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1309 _16309_/Q vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ _17901_/CLK _16917_/D vssd1 vssd1 vccd1 vccd1 _16917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17897_ _17897_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16848_ _18049_/CLK _16848_/D vssd1 vssd1 vccd1 vccd1 _16848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16779_ _18012_/CLK _16779_/D vssd1 vssd1 vccd1 vccd1 _16779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ hold2614/X _09325_/B _09319_/Y _14362_/A vssd1 vssd1 vccd1 vccd1 _09320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ hold944/X _16237_/Q _09273_/S vssd1 vssd1 vccd1 vccd1 hold945/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18449_ _18450_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08202_ hold1628/X _08213_/B _08201_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09182_ hold999/X _09230_/B vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _15705_/D sky130_fd_sc_hd__and2_1
XFILLER_0_172_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08064_ _15523_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3201 _18375_/Q vssd1 vssd1 vccd1 vccd1 hold3201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3212 _17421_/Q vssd1 vssd1 vccd1 vccd1 hold3212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3223 _14307_/X vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3234 _18023_/Q vssd1 vssd1 vccd1 vccd1 hold3234/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3245 _12956_/X vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2500 _15883_/Q vssd1 vssd1 vccd1 vccd1 hold2500/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3256 _17493_/Q vssd1 vssd1 vccd1 vccd1 hold3256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 _14095_/X vssd1 vssd1 vccd1 vccd1 _17850_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3267 _17489_/Q vssd1 vssd1 vccd1 vccd1 hold3267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 _15713_/Q vssd1 vssd1 vccd1 vccd1 hold2522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 _14669_/X vssd1 vssd1 vccd1 vccd1 _18125_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08966_ _12418_/A hold398/X vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__and2_1
XFILLER_0_228_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3278 _16337_/Q vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2544 _18299_/Q vssd1 vssd1 vccd1 vccd1 hold2544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3289 _17498_/Q vssd1 vssd1 vccd1 vccd1 hold3289/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2555 _15743_/Q vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_385_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1810 _14061_/X vssd1 vssd1 vccd1 vccd1 _17833_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2566 _18442_/Q vssd1 vssd1 vccd1 vccd1 hold2566/X sky130_fd_sc_hd__dlygate4sd3_1
X_07917_ hold2473/X _07918_/B _07916_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _07917_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1821 _17859_/Q vssd1 vssd1 vccd1 vccd1 hold1821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1832 _14833_/X vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2577 _18052_/Q vssd1 vssd1 vccd1 vccd1 hold2577/X sky130_fd_sc_hd__dlygate4sd3_1
X_08897_ _12386_/A hold455/X vssd1 vssd1 vccd1 vccd1 _16066_/D sky130_fd_sc_hd__and2_1
Xhold1843 _18198_/Q vssd1 vssd1 vccd1 vccd1 hold1843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 _15847_/Q vssd1 vssd1 vccd1 vccd1 hold2588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1854 _15232_/X vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2599 _15876_/Q vssd1 vssd1 vccd1 vccd1 hold2599/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_314_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17901_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1865 _18079_/Q vssd1 vssd1 vccd1 vccd1 hold1865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 _14899_/X vssd1 vssd1 vccd1 vccd1 _18235_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07848_ hold3021/X _07869_/B _07847_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _07848_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_233_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1887 _18223_/Q vssd1 vssd1 vccd1 vccd1 hold1887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1898 _09338_/X vssd1 vssd1 vccd1 vccd1 _16279_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09518_ hold2480/X _16330_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__mux2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ hold1511/X hold4295/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09449_ _09456_/D _09449_/B vssd1 vssd1 vccd1 vccd1 _16309_/D sky130_fd_sc_hd__nor2_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _17323_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ hold1783/X hold4325/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__mux2_1
X_12391_ hold17/X hold303/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ _15203_/A _14140_/B vssd1 vssd1 vccd1 vccd1 _14130_/X sky130_fd_sc_hd__or2_1
X_11342_ hold1454/X hold3924/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17505_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ hold1809/X _14094_/B _14060_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14061_/X
+ sky130_fd_sc_hd__o211a_1
X_11273_ hold1916/X hold4984/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5170 _16615_/Q vssd1 vssd1 vccd1 vccd1 hold5170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10224_ _10536_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ hold5983/X _13003_/Y _13011_/X _12531_/A vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5181 _10972_/X vssd1 vssd1 vccd1 vccd1 _16814_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5192 _16768_/Q vssd1 vssd1 vccd1 vccd1 hold5192/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4480 _13762_/X vssd1 vssd1 vccd1 vccd1 _17707_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17820_ _17883_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ _11103_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__or2_1
Xhold4491 _17026_/Q vssd1 vssd1 vccd1 vccd1 hold4491/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3790 _10144_/X vssd1 vssd1 vccd1 vccd1 _16538_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17751_ _18460_/CLK _17751_/D vssd1 vssd1 vccd1 vccd1 _17751_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ hold1702/X _14946_/B _14962_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14963_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ _10560_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _18182_/CLK _16702_/D vssd1 vssd1 vccd1 vccd1 _16702_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13914_ _15203_/A hold1531/X hold124/X vssd1 vssd1 vccd1 vccd1 _13915_/B sky130_fd_sc_hd__mux2_1
X_17682_ _17749_/CLK _17682_/D vssd1 vssd1 vccd1 vccd1 _17682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14894_ _14894_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14894_/X sky130_fd_sc_hd__or2_1
XFILLER_0_199_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16633_ _18221_/CLK _16633_/D vssd1 vssd1 vccd1 vccd1 _16633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13845_ hold3328/X _13779_/A _13844_/X vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16564_ _18152_/CLK _16564_/D vssd1 vssd1 vccd1 vccd1 _16564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13776_/X sky130_fd_sc_hd__or2_1
X_10988_ hold1263/X _16820_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10989_/B sky130_fd_sc_hd__mux2_1
X_18303_ _18303_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15515_ _15515_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ hold2662/X hold3197/X _12751_/S vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__mux2_1
X_16495_ _18374_/CLK _16495_/D vssd1 vssd1 vccd1 vccd1 _16495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ _18234_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15446_ _17320_/Q _09357_/A _09392_/A hold710/X vssd1 vssd1 vccd1 vccd1 _15446_/X
+ sky130_fd_sc_hd__a22o_1
X_12658_ hold2819/X _17397_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18165_ _18229_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
X_11609_ hold2508/X _17027_/Q _12365_/C vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__mux2_1
X_15377_ hold294/X _09357_/A _09386_/D _15895_/Q _15376_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12589_ hold905/X hold3230/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _17276_/CLK _17116_/D vssd1 vssd1 vccd1 vccd1 _17116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14328_ _14328_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__or2_1
X_18096_ _18212_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold406 hold406/A vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 hold417/A vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 hold428/A vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _17970_/CLK _17047_/D vssd1 vssd1 vccd1 vccd1 _17047_/Q sky130_fd_sc_hd__dfxtp_1
X_14259_ hold2974/X _14272_/B _14258_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _15121_/A vssd1 vssd1 vccd1 vccd1 _15555_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_221_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 hold972/X vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__buf_12
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ hold174/X hold195/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 input66/X vssd1 vssd1 vccd1 vccd1 hold1106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1117 _18261_/Q vssd1 vssd1 vccd1 vccd1 hold1117/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ hold98/X hold866/X _08779_/S vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__mux2_1
Xhold1128 _15803_/Q vssd1 vssd1 vccd1 vccd1 hold1128/X sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ _18305_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 _08461_/X vssd1 vssd1 vccd1 vccd1 _15859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08682_ _12444_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _15962_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _14984_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ _12696_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _16228_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09165_ hold2377/X _09164_/B _09164_/Y _12909_/A vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08116_ _14246_/A hold2118/X hold240/X vssd1 vssd1 vccd1 vccd1 _08117_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _15103_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08047_ hold752/X hold689/X hold764/X hold732/X vssd1 vssd1 vccd1 vccd1 _14627_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_226_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold940 hold940/A vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold951 hold951/A vssd1 vssd1 vccd1 vccd1 input2/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3020 _08412_/X vssd1 vssd1 vccd1 vccd1 _15836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3031 _18030_/Q vssd1 vssd1 vccd1 vccd1 hold3031/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3042 _14420_/X vssd1 vssd1 vccd1 vccd1 _18006_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3053 _18191_/Q vssd1 vssd1 vccd1 vccd1 hold3053/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3064 _14639_/X vssd1 vssd1 vccd1 vccd1 _18110_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09998_ _16490_/Q _11159_/B _11159_/C vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__and3_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3075 _18134_/Q vssd1 vssd1 vccd1 vccd1 hold3075/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2330 _14177_/X vssd1 vssd1 vccd1 vccd1 _17889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3086 _18167_/Q vssd1 vssd1 vccd1 vccd1 hold3086/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2341 _18128_/Q vssd1 vssd1 vccd1 vccd1 hold2341/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3097 _18115_/Q vssd1 vssd1 vccd1 vccd1 hold3097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 _14267_/X vssd1 vssd1 vccd1 vccd1 _17932_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08949_ hold596/X hold876/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold877/A sky130_fd_sc_hd__mux2_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2363 _15581_/Q vssd1 vssd1 vccd1 vccd1 hold2363/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2374 _08304_/X vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _18042_/Q vssd1 vssd1 vccd1 vccd1 hold1640/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2385 _08097_/X vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2396 _09159_/X vssd1 vssd1 vccd1 vccd1 _16192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 _14121_/X vssd1 vssd1 vccd1 vccd1 _17862_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1662 _15757_/Q vssd1 vssd1 vccd1 vccd1 hold1662/X sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ hold2612/X hold4543/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__mux2_1
Xhold1673 _14929_/X vssd1 vssd1 vccd1 vccd1 _18249_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1684 _15620_/Q vssd1 vssd1 vccd1 vccd1 hold1684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1695 _18252_/Q vssd1 vssd1 vccd1 vccd1 hold1695/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _11694_/A _10911_/B vssd1 vssd1 vccd1 vccd1 _10911_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ hold2522/X hold3736/X _13877_/C vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__mux2_1
X_13630_ hold5713/X _13829_/B _13629_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13630_/X
+ sky130_fd_sc_hd__o211a_1
X_10842_ _11121_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ hold3531/X _13847_/B _13560_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ _11064_/A _10773_/B vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ hold230/X _15486_/A2 _09357_/B hold409/X vssd1 vssd1 vccd1 vccd1 _15300_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12512_ _09342_/A hold2124/X _07802_/Y _12511_/X vssd1 vssd1 vccd1 vccd1 _12512_/X
+ sky130_fd_sc_hd__o211a_1
X_16280_ _18460_/CLK _16280_/D vssd1 vssd1 vccd1 vccd1 _16280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13492_ hold3482/X _13886_/B _13491_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15231_ _15231_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__or2_1
X_12443_ hold150/X hold415/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold416/A sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ hold1204/X _15165_/B _15161_/Y _15162_/C1 vssd1 vssd1 vccd1 vccd1 _15162_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _17282_/Q _12374_/B _13556_/S vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14113_ hold1446/X _14142_/B _14112_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _12213_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__or2_1
X_15093_ _15201_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14044_ _14330_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14044_/X sky130_fd_sc_hd__or2_1
X_11256_ _11553_/A _11256_/B vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_236_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18153_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_235_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ hold4944/X _10649_/B _10206_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10207_/X
+ sky130_fd_sc_hd__o211a_1
X_11187_ hold4632/X _11103_/A _11186_/X vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10138_ hold3839/X _11198_/B _10137_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _10138_/X
+ sky130_fd_sc_hd__o211a_1
X_17803_ _17890_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _18415_/CLK _15995_/D vssd1 vssd1 vccd1 vccd1 _15995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _17734_/CLK _17734_/D vssd1 vssd1 vccd1 vccd1 _17734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ _10603_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _16513_/D sky130_fd_sc_hd__nor2_1
X_14946_ _14946_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17665_ _17695_/CLK _17665_/D vssd1 vssd1 vccd1 vccd1 _17665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14877_ hold1174/X _14880_/B _14876_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14877_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16616_ _18210_/CLK _16616_/D vssd1 vssd1 vccd1 vccd1 _16616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ _13864_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _17729_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17596_ _17723_/CLK _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16547_ _18216_/CLK _16547_/D vssd1 vssd1 vccd1 vccd1 _16547_/Q sky130_fd_sc_hd__dfxtp_1
X_13759_ hold4147/X _13886_/B _13758_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16478_ _18383_/CLK _16478_/D vssd1 vssd1 vccd1 vccd1 _16478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18217_ _18219_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15429_ hold769/X _09386_/A _15427_/X vssd1 vssd1 vccd1 vccd1 _15432_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_182_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18148_ _18186_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5906 _07797_/X vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5917 _16911_/Q vssd1 vssd1 vccd1 vccd1 hold5917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5928 _17547_/Q vssd1 vssd1 vccd1 vccd1 hold5928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__clkbuf_8
Xhold214 input27/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5939 _17554_/Q vssd1 vssd1 vccd1 vccd1 hold5939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _18143_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold236 hold729/X vssd1 vssd1 vccd1 vccd1 hold730/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold28/X vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _09963_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__or2_1
Xfanout705 _12396_/A vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout716 _13037_/A vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__clkbuf_4
X_09852_ _09936_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__or2_1
Xfanout727 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__clkbuf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout738 _15473_/A vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__buf_4
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _08377_/A vssd1 vssd1 vccd1 vccd1 _08111_/A sky130_fd_sc_hd__clkbuf_4
X_08803_ _08868_/B _12380_/B _13046_/D vssd1 vssd1 vccd1 vccd1 _08808_/S sky130_fd_sc_hd__or3_2
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10191_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08734_ _12418_/A hold855/X vssd1 vssd1 vccd1 vccd1 _15987_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ hold554/X hold641/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold642/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _13043_/C hold990/X vssd1 vssd1 vccd1 vccd1 _13034_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ hold2579/X _09218_/B _09216_/Y _12912_/A vssd1 vssd1 vccd1 vccd1 _09217_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09148_ _15531_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ hold1063/X _09119_/A2 _09078_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11110_ hold5565/X _11753_/B _11109_/X _14538_/C1 vssd1 vssd1 vccd1 vccd1 _11110_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _12273_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold781 hold781/A vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold792 hold792/A vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ hold5583/X _11156_/B _11040_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _11041_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _17899_/Q vssd1 vssd1 vccd1 vccd1 hold2160/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2171 _14663_/X vssd1 vssd1 vccd1 vccd1 _18122_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _15193_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__or2_1
XFILLER_0_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 _15565_/Q vssd1 vssd1 vccd1 vccd1 hold2182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_232_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _17736_/CLK _15780_/D vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_235_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2193 _08004_/X vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ hold3273/X _12991_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_231_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1470 _18393_/Q vssd1 vssd1 vccd1 vccd1 hold1470/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ hold1529/X _14714_/B _14730_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14731_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1481 _18379_/Q vssd1 vssd1 vccd1 vccd1 hold1481/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1492 _14945_/X vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _12267_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17450_ _17878_/CLK _17450_/D vssd1 vssd1 vccd1 vccd1 _17450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14878_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14662_/Y sky130_fd_sc_hd__nand2_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ _13794_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__or2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _18386_/CLK _16401_/D vssd1 vssd1 vccd1 vccd1 _16401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13613_ hold2727/X hold4166/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17485_/CLK _17381_/D vssd1 vssd1 vccd1 vccd1 _17381_/Q sky130_fd_sc_hd__dfxtp_1
X_10825_ hold5467/X _11207_/B _10824_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10825_/X
+ sky130_fd_sc_hd__o211a_1
X_14593_ hold3189/X _14610_/B _14592_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16332_ _18309_/CLK _16332_/D vssd1 vssd1 vccd1 vccd1 _16332_/Q sky130_fd_sc_hd__dfxtp_1
X_13544_ _15820_/Q _17635_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ hold4279/X _11729_/B _10755_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _10756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16263_ _17365_/CLK _16263_/D vssd1 vssd1 vccd1 vccd1 _16263_/Q sky130_fd_sc_hd__dfxtp_1
X_13475_ hold1145/X _17612_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ hold5196/X _11738_/B _10686_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _10687_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18002_ _18035_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ hold1565/X _15221_/B _15213_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15214_/X
+ sky130_fd_sc_hd__o211a_1
X_12426_ _12426_/A hold861/X vssd1 vssd1 vccd1 vccd1 _17306_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16194_ _17478_/CLK _16194_/D vssd1 vssd1 vccd1 vccd1 _16194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_417_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17260_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15145_ _15199_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12357_ hold4779/X _12261_/A _12356_/X vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ hold5256/X _12329_/B _11307_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11308_/X
+ sky130_fd_sc_hd__o211a_1
X_15076_ hold1787/X _15111_/B _15075_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15076_/X
+ sky130_fd_sc_hd__o211a_1
X_12288_ _12288_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__or2_1
X_14027_ hold2939/X _14040_/B _14026_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14027_/X
+ sky130_fd_sc_hd__o211a_1
X_11239_ hold5014/X _12299_/B _11238_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _11239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15978_ _17297_/CLK _15978_/D vssd1 vssd1 vccd1 vccd1 hold633/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ hold1672/X _14952_/B _14928_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _14929_/X
+ sky130_fd_sc_hd__o211a_1
X_17717_ _17749_/CLK _17717_/D vssd1 vssd1 vccd1 vccd1 _17717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08450_ _15509_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08450_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17648_ _17739_/CLK _17648_/D vssd1 vssd1 vccd1 vccd1 _17648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _15822_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17579_ _17736_/CLK _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ hold312/X hold372/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold373/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5703 _17666_/Q vssd1 vssd1 vccd1 vccd1 hold5703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5714 _13630_/X vssd1 vssd1 vccd1 vccd1 _17663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_158_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18237_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5725 _17654_/Q vssd1 vssd1 vccd1 vccd1 hold5725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5736 _13354_/X vssd1 vssd1 vccd1 vccd1 _17571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5747 _17664_/Q vssd1 vssd1 vccd1 vccd1 hold5747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5758 _13387_/X vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5769 hold5925/X vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout502 _10400_/S vssd1 vssd1 vccd1 vccd1 _11093_/S sky130_fd_sc_hd__buf_4
X_09904_ hold5252/X _11159_/B _09903_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09904_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout513 _10589_/C vssd1 vssd1 vccd1 vccd1 _10649_/C sky130_fd_sc_hd__clkbuf_8
Xfanout524 _09285_/Y vssd1 vssd1 vccd1 vccd1 _09338_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout535 _09066_/Y vssd1 vssd1 vccd1 vccd1 _09106_/B sky130_fd_sc_hd__buf_4
Xfanout546 hold205/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__buf_6
X_09835_ hold3827/X _10019_/B _09834_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09835_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout557 hold239/X vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__buf_4
Xfanout568 _07916_/B vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__buf_8
Xfanout579 _13057_/X vssd1 vssd1 vccd1 vccd1 _13250_/S sky130_fd_sc_hd__buf_8
XFILLER_0_214_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09766_ hold3992/X _10034_/B _09765_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_240_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ hold210/X hold816/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold817/A sky130_fd_sc_hd__mux2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ hold3381/X _10025_/B _09696_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _09697_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08648_ _12408_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _15946_/D sky130_fd_sc_hd__and2_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08579_ _15414_/A hold319/X vssd1 vssd1 vccd1 vccd1 _15913_/D sky130_fd_sc_hd__and2_1
XFILLER_0_37_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10610_ _16694_/Q _10646_/B _10997_/S vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__and3_1
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ hold5230/X _12314_/B _11589_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11590_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ hold1970/X hold4986/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13260_ hold4962/X _13259_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__mux2_2
X_10472_ hold1831/X _16648_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ hold5022/X _12308_/B _12210_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _12211_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13191_ _13199_/A1 _13189_/X _13190_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ hold4187/X _13868_/B _12141_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _12142_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12073_ hold3450/X _12347_/B _12072_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _12073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16950_ _17935_/CLK _16950_/D vssd1 vssd1 vccd1 vccd1 _16950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15901_ _17304_/CLK _15901_/D vssd1 vssd1 vccd1 vccd1 hold801/A sky130_fd_sc_hd__dfxtp_1
X_11024_ hold1823/X hold5020/X _11216_/C vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__mux2_1
X_16881_ _18050_/CLK _16881_/D vssd1 vssd1 vccd1 vccd1 _16881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15832_ _17721_/CLK _15832_/D vssd1 vssd1 vccd1 vccd1 _15832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _17749_/CLK _15763_/D vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__and2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _15215_/A _14714_/B vssd1 vssd1 vccd1 vccd1 _14714_/Y sky130_fd_sc_hd__nand2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17879_/CLK _17502_/D vssd1 vssd1 vccd1 vccd1 _17502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ hold5100/X _13798_/A2 _11925_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15694_ _17166_/CLK _15694_/D vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17433_ _18453_/CLK _17433_/D vssd1 vssd1 vccd1 vccd1 _17433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ hold3093/X _14664_/B _14644_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14645_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11857_ hold4317/X _12374_/B _11856_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _11857_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10808_ hold2477/X _16760_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
X_17364_ _17365_/CLK _17364_/D vssd1 vssd1 vccd1 vccd1 _17364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ _15131_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__or2_1
X_11788_ _12340_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _17086_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_138_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16315_ _16323_/CLK _16315_/D vssd1 vssd1 vccd1 vccd1 _16315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13527_ _13623_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17295_ _17298_/CLK _17295_/D vssd1 vssd1 vccd1 vccd1 hold868/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ hold2759/X hold3850/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16246_ _17425_/CLK hold183/X vssd1 vssd1 vccd1 vccd1 _16246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13458_ _13746_/A _13458_/B vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_251_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ hold118/X hold803/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_140_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16177_ _17482_/CLK _16177_/D vssd1 vssd1 vccd1 vccd1 _16177_/Q sky130_fd_sc_hd__dfxtp_1
X_13389_ _13773_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 _17524_/Q vssd1 vssd1 vccd1 vccd1 io_out sky130_fd_sc_hd__buf_12
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4309 _17701_/Q vssd1 vssd1 vccd1 vccd1 hold4309/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput116 hold5874/X vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_12
Xoutput127 hold5844/X vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_12
X_15128_ _15128_/A hold393/X vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__or2_4
Xoutput138 hold5877/X vssd1 vssd1 vccd1 vccd1 hold5878/A sky130_fd_sc_hd__buf_6
XFILLER_0_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3608 _10647_/Y vssd1 vssd1 vccd1 vccd1 _10648_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3619 _16375_/Q vssd1 vssd1 vccd1 vccd1 hold3619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15059_ hold367/X hold844/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold845/A sky130_fd_sc_hd__mux2_1
X_07950_ _14854_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_220_1359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2907 _17888_/Q vssd1 vssd1 vccd1 vccd1 hold2907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 _14474_/X vssd1 vssd1 vccd1 vccd1 _18032_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2929 _15599_/Q vssd1 vssd1 vccd1 vccd1 hold2929/X sky130_fd_sc_hd__dlygate4sd3_1
X_07881_ _15559_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_218_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09620_ hold1283/X hold3808/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_207_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ hold1695/X _13198_/A _10055_/C vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_222_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08502_ hold752/X hold732/X hold764/X hold689/X vssd1 vssd1 vccd1 vccd1 _14897_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09482_ hold895/X _09482_/B vssd1 vssd1 vccd1 vccd1 _09484_/C sky130_fd_sc_hd__or2_1
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ _14774_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08364_ _15533_/A hold2523/X hold134/X vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_339_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17280_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ _14854_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5500 _13384_/X vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5511 _17270_/Q vssd1 vssd1 vccd1 vccd1 hold5511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5522 _10984_/X vssd1 vssd1 vccd1 vccd1 _16818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5533 _17081_/Q vssd1 vssd1 vccd1 vccd1 hold5533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5544 _10945_/X vssd1 vssd1 vccd1 vccd1 _16805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4810 _09550_/X vssd1 vssd1 vccd1 vccd1 _16340_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5555 _16948_/Q vssd1 vssd1 vccd1 vccd1 hold5555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4821 _16506_/Q vssd1 vssd1 vccd1 vccd1 hold4821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5566 _11110_/X vssd1 vssd1 vccd1 vccd1 _16860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4832 _09943_/X vssd1 vssd1 vccd1 vccd1 _16471_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5577 _17075_/Q vssd1 vssd1 vccd1 vccd1 hold5577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4843 _16410_/Q vssd1 vssd1 vccd1 vccd1 hold4843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5588 _11386_/X vssd1 vssd1 vccd1 vccd1 _16952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4854 _10438_/X vssd1 vssd1 vccd1 vccd1 _16636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5599 _17206_/Q vssd1 vssd1 vccd1 vccd1 hold5599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4865 _16579_/Q vssd1 vssd1 vccd1 vccd1 hold4865/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4876 _10387_/X vssd1 vssd1 vccd1 vccd1 _16619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout310 _10467_/A vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__buf_4
Xfanout321 _10470_/A vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__buf_4
Xhold4887 _16760_/Q vssd1 vssd1 vccd1 vccd1 hold4887/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout332 _09564_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__clkbuf_4
Xhold4898 _10177_/X vssd1 vssd1 vccd1 vccd1 _16549_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout343 _09056_/S vssd1 vssd1 vccd1 vccd1 _09062_/S sky130_fd_sc_hd__buf_8
Xfanout354 _08627_/S vssd1 vssd1 vccd1 vccd1 _08655_/S sky130_fd_sc_hd__buf_8
Xfanout365 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15165_/B sky130_fd_sc_hd__clkbuf_8
Xfanout376 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__buf_6
XFILLER_0_214_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09818_ _18341_/Q _16430_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__mux2_1
Xfanout387 _14680_/Y vssd1 vssd1 vccd1 vccd1 _14720_/B sky130_fd_sc_hd__buf_8
Xfanout398 _14411_/B vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__buf_6
XFILLER_0_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17985_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09749_ _18318_/Q _16407_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12760_ hold2752/X _17431_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__mux2_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ hold1505/X hold3784/X _11711_/S vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ hold1422/X hold3785/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ hold2066/X _14433_/B _14429_/Y _12981_/A vssd1 vssd1 vccd1 vccd1 _14430_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ hold1545/X _17038_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ _14988_/A hold2966/X hold333/X vssd1 vssd1 vccd1 vccd1 _14362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ hold2274/X hold5647/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 input18/A vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_6
X_16100_ _18418_/CLK _16100_/D vssd1 vssd1 vccd1 vccd1 hold397/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _13305_/X _13311_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_135_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_6
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or2_1
X_17080_ _17894_/CLK _17080_/D vssd1 vssd1 vccd1 vccd1 _17080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14292_ _14972_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14292_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_18_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_18_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_16031_ _18401_/CLK _16031_/D vssd1 vssd1 vccd1 vccd1 hold768/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13243_ _13242_/X _16923_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__mux2_2
X_10455_ _10998_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ _13174_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ _10482_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12125_ hold2717/X hold4201/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_209_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17982_ _18014_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12056_ hold1785/X _17176_/Q _12344_/C vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__mux2_1
X_16933_ _17875_/CLK _16933_/D vssd1 vssd1 vccd1 vccd1 _16933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11103_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__or2_1
X_16864_ _18065_/CLK _16864_/D vssd1 vssd1 vccd1 vccd1 _16864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15815_ _17666_/CLK _15815_/D vssd1 vssd1 vccd1 vccd1 _15815_/Q sky130_fd_sc_hd__dfxtp_1
X_16795_ _17996_/CLK _16795_/D vssd1 vssd1 vccd1 vccd1 _16795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15746_ _17747_/CLK _15746_/D vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12958_ hold2455/X _17497_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ hold2616/X _17127_/Q _12302_/C vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _17265_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ hold2923/X _17474_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_57_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_57_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14628_ _14968_/A _14676_/B vssd1 vssd1 vccd1 vccd1 _14628_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17416_ _17429_/CLK _17416_/D vssd1 vssd1 vccd1 vccd1 _17416_/Q sky130_fd_sc_hd__dfxtp_1
X_18396_ _18396_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _17347_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _17347_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_432_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17677_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14559_ _14968_/A _14557_/Y hold1219/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14559_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _15539_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08080_/X sky130_fd_sc_hd__or2_1
X_17278_ _17278_/CLK _17278_/D vssd1 vssd1 vccd1 vccd1 _17278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16229_ _17431_/CLK _16229_/D vssd1 vssd1 vccd1 vccd1 _16229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4106 _10735_/X vssd1 vssd1 vccd1 vccd1 _16735_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4117 hold5891/X vssd1 vssd1 vccd1 vccd1 hold5892/A sky130_fd_sc_hd__buf_6
XFILLER_0_109_1388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4128 _12238_/X vssd1 vssd1 vccd1 vccd1 _17236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4139 _17406_/Q vssd1 vssd1 vccd1 vccd1 hold4139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3405 _16397_/Q vssd1 vssd1 vccd1 vccd1 hold3405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3416 _12617_/X vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08982_ _12436_/A hold297/X vssd1 vssd1 vccd1 vccd1 _16108_/D sky130_fd_sc_hd__and2_1
Xhold3427 _09529_/X vssd1 vssd1 vccd1 vccd1 _16333_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3438 _16710_/Q vssd1 vssd1 vccd1 vccd1 hold3438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2704 _14585_/X vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3449 _12253_/X vssd1 vssd1 vccd1 vccd1 _17241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2715 _15830_/Q vssd1 vssd1 vccd1 vccd1 hold2715/X sky130_fd_sc_hd__dlygate4sd3_1
X_07933_ hold2590/X _07924_/B _07932_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _07933_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2726 _14087_/X vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2737 _17898_/Q vssd1 vssd1 vccd1 vccd1 hold2737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2748 _16217_/Q vssd1 vssd1 vccd1 vccd1 hold2748/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2759 _17938_/Q vssd1 vssd1 vccd1 vccd1 hold2759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07864_ hold2212/X _07869_/B _07863_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 _07864_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09603_ _09987_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07795_ _18459_/Q hold1412/X _09342_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _07795_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_218_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _09933_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09472_/D _09465_/B vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__nor2_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08416_ hold2867/X _08440_/A2 _08415_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _09386_/B _09369_/B _18458_/Q vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_173_wb_clk_i clkbuf_6_48_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18351_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08347_ _08391_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__and2_1
XFILLER_0_188_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08278_ _15557_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6020 data_in[3] vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6031 _18402_/Q vssd1 vssd1 vccd1 vccd1 hold6031/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6042 _16518_/Q vssd1 vssd1 vccd1 vccd1 hold6042/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5330 _16633_/Q vssd1 vssd1 vccd1 vccd1 hold5330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10240_ hold4899/X _10649_/B _10239_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10240_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5341 _12226_/X vssd1 vssd1 vccd1 vccd1 _17232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5352 _16976_/Q vssd1 vssd1 vccd1 vccd1 hold5352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5363 _09712_/X vssd1 vssd1 vccd1 vccd1 _16394_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5374 _10300_/X vssd1 vssd1 vccd1 vccd1 _16590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4640 _10632_/Y vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5385 _16957_/Q vssd1 vssd1 vccd1 vccd1 hold5385/X sky130_fd_sc_hd__dlygate4sd3_1
X_10171_ hold4865/X _10649_/B _10170_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10171_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4651 _16336_/Q vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5396 _11254_/X vssd1 vssd1 vccd1 vccd1 _16908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4662 _16924_/Q vssd1 vssd1 vccd1 vccd1 hold4662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4673 _12300_/Y vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4684 _11718_/Y vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3950 _16631_/Q vssd1 vssd1 vccd1 vccd1 hold3950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4695 _17107_/Q vssd1 vssd1 vccd1 vccd1 hold4695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3961 _09532_/X vssd1 vssd1 vccd1 vccd1 _16334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3972 _16627_/Q vssd1 vssd1 vccd1 vccd1 hold3972/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout151 _12827_/S vssd1 vssd1 vccd1 vccd1 _12809_/S sky130_fd_sc_hd__buf_6
Xhold3983 _10450_/X vssd1 vssd1 vccd1 vccd1 _16640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout162 _12293_/B vssd1 vssd1 vccd1 vccd1 _13811_/B sky130_fd_sc_hd__buf_4
XFILLER_0_233_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3994 _17240_/Q vssd1 vssd1 vccd1 vccd1 hold3994/X sky130_fd_sc_hd__dlygate4sd3_1
X_13930_ hold181/A _17771_/Q hold124/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__mux2_1
Xfanout173 _11617_/A2 vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__clkbuf_8
Xfanout184 _13777_/A2 vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout195 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _12274_/A2 sky130_fd_sc_hd__buf_4
X_13861_ _13888_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _17740_/D sky130_fd_sc_hd__nor2_1
X_15600_ _17283_/CLK _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12812_ hold3183/X _12811_/X _12827_/S vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16580_ _18232_/CLK _16580_/D vssd1 vssd1 vccd1 vccd1 _16580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13792_ hold4405/X _13880_/B _13791_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15531_ _15531_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__or2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ hold3205/X _12742_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18316_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15480_/A _15462_/B _15462_/C _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_166_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12674_ hold3847/X _12673_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17266_/CLK _17201_/D vssd1 vssd1 vccd1 vccd1 _17201_/Q sky130_fd_sc_hd__dfxtp_1
X_14413_ _15201_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__or2_1
X_18181_ _18181_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _12204_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15393_ _15481_/A1 _15385_/X _15392_/X _15481_/B1 _18413_/Q vssd1 vssd1 vccd1 vccd1
+ _15393_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_155_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17132_ _17260_/CLK _17132_/D vssd1 vssd1 vccd1 vccd1 _17132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_231_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14344_ _14344_/A _14344_/B vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__and2_1
XFILLER_0_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11556_ _12219_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or2_1
X_10507_ _10601_/A _10619_/B _10506_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _10507_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17063_ _18427_/CLK _17063_/D vssd1 vssd1 vccd1 vccd1 _17063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14275_ hold2512/X _14272_/B _14274_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14275_/X
+ sky130_fd_sc_hd__o211a_1
X_11487_ _12243_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__or2_1
X_16014_ _18421_/CLK _16014_/D vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13226_ _17579_/Q _17113_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ hold4853/X _10625_/B _10437_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13157_ _13156_/X hold3547/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ hold4028/X _10565_/B _10368_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12204_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13081_/X _13087_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17529_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_178_1342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17997_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12039_ _12231_/A _12039_/B vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__or2_1
X_16916_ _17858_/CLK _16916_/D vssd1 vssd1 vccd1 vccd1 _16916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17896_ _17896_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16847_ _17952_/CLK _16847_/D vssd1 vssd1 vccd1 vccd1 _16847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16778_ _18043_/CLK _16778_/D vssd1 vssd1 vccd1 vccd1 _16778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15729_ _17700_/CLK _15729_/D vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_6_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09250_ _12759_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _16236_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _18448_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08201_ _14529_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ hold1181/X _09218_/B _09180_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__o211a_1
X_18379_ _18379_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08132_ _15537_/A hold2438/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ hold2227/X _08097_/A2 _08062_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _08063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3202 _15190_/X vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3213 _18055_/Q vssd1 vssd1 vccd1 vccd1 hold3213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3224 _17467_/Q vssd1 vssd1 vccd1 vccd1 hold3224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3235 _14456_/X vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3246 _16329_/Q vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2501 _08512_/X vssd1 vssd1 vccd1 vccd1 _15883_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08965_ hold346/X hold397/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold398/A sky130_fd_sc_hd__mux2_1
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3257 _17357_/Q vssd1 vssd1 vccd1 vccd1 hold3257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 _17936_/Q vssd1 vssd1 vccd1 vccd1 hold2512/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3268 _12938_/X vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _15814_/Q vssd1 vssd1 vccd1 vccd1 hold2523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3279 _10020_/Y vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 _15694_/Q vssd1 vssd1 vccd1 vccd1 hold2534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 _14919_/X vssd1 vssd1 vccd1 vccd1 _18244_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2545 _17983_/Q vssd1 vssd1 vccd1 vccd1 hold2545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 _18372_/Q vssd1 vssd1 vccd1 vccd1 hold1811/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2556 _08214_/X vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07916_ _15539_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07916_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1822 _14115_/X vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08896_ hold454/X _16066_/Q _08928_/S vssd1 vssd1 vccd1 vccd1 hold455/A sky130_fd_sc_hd__mux2_1
Xhold2567 _15532_/X vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 _16323_/Q vssd1 vssd1 vccd1 vccd1 hold1833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 _14516_/X vssd1 vssd1 vccd1 vccd1 _18052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _14821_/X vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 _08434_/X vssd1 vssd1 vccd1 vccd1 _15847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1855 _18107_/Q vssd1 vssd1 vccd1 vccd1 hold1855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 _14575_/X vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07847_ _15525_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07847_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1877 _16278_/Q vssd1 vssd1 vccd1 vccd1 hold1877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1888 _14873_/X vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1899 _18081_/Q vssd1 vssd1 vccd1 vccd1 hold1899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09517_ hold3361/X _10013_/B _09516_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09517_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_354_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17612_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09448_ _09447_/A _09444_/X _09484_/B vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__o21ai_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ _17326_/Q _09357_/A _09392_/C hold504/X _09378_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_81_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11410_ hold5603/X _12365_/B _11409_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _12416_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _17288_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ hold3910/X _11726_/B _11340_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11341_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _14972_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ hold5509/X _11753_/B _11271_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11272_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5160 _17157_/Q vssd1 vssd1 vccd1 vccd1 hold5160/X sky130_fd_sc_hd__dlygate4sd3_1
X_13011_ _14974_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__or2_1
X_10223_ hold2407/X _16565_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__mux2_1
Xhold5171 _10279_/X vssd1 vssd1 vccd1 vccd1 _16583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5182 _16648_/Q vssd1 vssd1 vccd1 vccd1 hold5182/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5193 _10738_/X vssd1 vssd1 vccd1 vccd1 _16736_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4470 _11596_/X vssd1 vssd1 vccd1 vccd1 _17022_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ hold2447/X hold4619/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__mux2_1
Xhold4481 _16400_/Q vssd1 vssd1 vccd1 vccd1 hold4481/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4492 _11512_/X vssd1 vssd1 vccd1 vccd1 _16994_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3780 _12704_/X vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14962_ _15231_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14962_/X sky130_fd_sc_hd__or2_1
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ _18460_/CLK _17750_/D vssd1 vssd1 vccd1 vccd1 _17750_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3791 _17584_/Q vssd1 vssd1 vccd1 vccd1 hold3791/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ hold2087/X hold3543/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__mux2_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _18225_/CLK _16701_/D vssd1 vssd1 vccd1 vccd1 _16701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ _13923_/A _13913_/B vssd1 vssd1 vccd1 vccd1 _17762_/D sky130_fd_sc_hd__and2_1
X_14893_ hold1739/X _14880_/B _14892_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _14893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17681_ _17681_/CLK _17681_/D vssd1 vssd1 vccd1 vccd1 _17681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16632_ _17968_/CLK _16632_/D vssd1 vssd1 vccd1 vccd1 _16632_/Q sky130_fd_sc_hd__dfxtp_1
X_13844_ _17735_/Q _13883_/B _13874_/C vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__and3_1
XFILLER_0_199_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16563_ _18175_/CLK _16563_/D vssd1 vssd1 vccd1 vccd1 _16563_/Q sky130_fd_sc_hd__dfxtp_1
X_13775_ hold2051/X _17712_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ hold4703/X _11177_/B _10986_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10987_/X
+ sky130_fd_sc_hd__o211a_1
X_18302_ _18421_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _12738_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _17418_/D sky130_fd_sc_hd__and2_1
X_15514_ hold2054/X _15507_/Y _15513_/X _12780_/A vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__o211a_1
X_16494_ _18342_/CLK _16494_/D vssd1 vssd1 vccd1 vccd1 _16494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ hold316/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__or2_1
X_18233_ _18233_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12657_ _12657_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _17395_/D sky130_fd_sc_hd__and2_1
XFILLER_0_210_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ hold4549/X _12344_/B _11607_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _11608_/X
+ sky130_fd_sc_hd__o211a_1
X_15376_ _17341_/Q _15479_/B1 _09362_/D hold372/X vssd1 vssd1 vccd1 vccd1 _15376_/X
+ sky130_fd_sc_hd__a22o_1
X_18164_ _18164_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ _14362_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _17372_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14327_ hold2477/X _14326_/B _14326_/Y _14392_/A vssd1 vssd1 vccd1 vccd1 _14327_/X
+ sky130_fd_sc_hd__o211a_1
X_17115_ _17261_/CLK _17115_/D vssd1 vssd1 vccd1 vccd1 _17115_/Q sky130_fd_sc_hd__dfxtp_1
X_18095_ _18141_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ hold4227/X _11729_/B _11538_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 hold407/A vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17046_ _17935_/CLK _17046_/D vssd1 vssd1 vccd1 vccd1 _17046_/Q sky130_fd_sc_hd__dfxtp_1
Xhold429 hold429/A vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ _15099_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _13209_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ hold1448/X _14202_/B _14188_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14189_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout909 _15121_/A vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__buf_4
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08750_ _15264_/A hold164/X vssd1 vssd1 vccd1 vccd1 _15995_/D sky130_fd_sc_hd__and2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 hold1107/A vssd1 vssd1 vccd1 vccd1 hold1107/X sky130_fd_sc_hd__clkbuf_8
Xhold1118 _14953_/X vssd1 vssd1 vccd1 vccd1 _18261_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _18044_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _17989_/Q vssd1 vssd1 vccd1 vccd1 hold1129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08681_ hold174/X hold363/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__mux2_1
X_17879_ _17879_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09302_ hold1547/X _09338_/A2 _09301_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09302_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _15509_/A hold1422/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ _15547_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ hold1775/X _09106_/B _09094_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08046_ hold1785/X _08033_/B _08045_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _08046_/X
+ sky130_fd_sc_hd__o211a_1
Xhold930 hold930/A vssd1 vssd1 vccd1 vccd1 hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 hold941/A vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold952 input2/X vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold974 hold974/A vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3010 _18009_/Q vssd1 vssd1 vccd1 vccd1 hold3010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 input48/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 _15569_/Q vssd1 vssd1 vccd1 vccd1 hold3021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 _14470_/X vssd1 vssd1 vccd1 vccd1 _18030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3043 _18146_/Q vssd1 vssd1 vccd1 vccd1 hold3043/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3054 _14807_/X vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _11203_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _16489_/D sky130_fd_sc_hd__nor2_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3065 _16163_/Q vssd1 vssd1 vccd1 vccd1 hold3065/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2320 _13981_/X vssd1 vssd1 vccd1 vccd1 _17795_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2331 _17785_/Q vssd1 vssd1 vccd1 vccd1 hold2331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3076 _14689_/X vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3087 _14757_/X vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2342 _14675_/X vssd1 vssd1 vccd1 vccd1 _18128_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08948_ _12412_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _16091_/D sky130_fd_sc_hd__and2_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3098 _14649_/X vssd1 vssd1 vccd1 vccd1 _18115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2353 _18180_/Q vssd1 vssd1 vccd1 vccd1 hold2353/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 _07872_/X vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2375 _15759_/Q vssd1 vssd1 vccd1 vccd1 hold2375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 _15861_/Q vssd1 vssd1 vccd1 vccd1 hold1630/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _14494_/X vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _15706_/Q vssd1 vssd1 vccd1 vccd1 hold2386/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2397 _18085_/Q vssd1 vssd1 vccd1 vccd1 hold2397/X sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ _15414_/A hold89/X vssd1 vssd1 vccd1 vccd1 _16057_/D sky130_fd_sc_hd__and2_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1652 _15841_/Q vssd1 vssd1 vccd1 vccd1 hold1652/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1663 _08245_/X vssd1 vssd1 vccd1 vccd1 _15757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _15752_/Q vssd1 vssd1 vccd1 vccd1 hold1674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ hold1393/X hold4419/X _11768_/C vssd1 vssd1 vccd1 vccd1 _10911_/B sky130_fd_sc_hd__mux2_1
Xhold1685 _07955_/X vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1696 _14935_/X vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ hold4340/X _12274_/A2 _11889_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ hold2112/X hold5573/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_212_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _13746_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10772_ hold1365/X hold5300/X _11159_/C vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _07809_/X _12510_/Y _13048_/A hold2124/X vssd1 vssd1 vccd1 vccd1 _12511_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_13491_ _13779_/A _13491_/B vssd1 vssd1 vccd1 vccd1 _13491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ hold2695/X _15221_/B _15229_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15230_/X
+ sky130_fd_sc_hd__o211a_1
X_12442_ _15364_/A hold772/X vssd1 vssd1 vccd1 vccd1 _17314_/D sky130_fd_sc_hd__and2_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15161_ _15215_/A _15165_/B vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _13888_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _17281_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_62_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ hold915/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11324_ hold1525/X hold3829/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__mux2_1
X_15092_ hold1985/X _15111_/B _15091_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _15092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14043_ hold2258/X _14038_/B _14042_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14043_/X
+ sky130_fd_sc_hd__o211a_1
X_11255_ hold2642/X hold4674/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11256_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10554_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__or2_1
XTAP_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _16886_/Q _11198_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__and3_1
XTAP_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17802_ _17834_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ _10830_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__or2_1
XTAP_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _18407_/CLK _15994_/D vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_276_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18234_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17733_ _17739_/CLK _17733_/D vssd1 vssd1 vccd1 vccd1 _17733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10068_ _13294_/A _10560_/A _10067_/X vssd1 vssd1 vccd1 vccd1 _10068_/Y sky130_fd_sc_hd__a21oi_1
X_14945_ hold1491/X _14946_/B _14944_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_205_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18382_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_215_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17664_ _17696_/CLK _17664_/D vssd1 vssd1 vccd1 vccd1 _17664_/Q sky130_fd_sc_hd__dfxtp_1
X_14876_ _15215_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16615_ _18205_/CLK _16615_/D vssd1 vssd1 vccd1 vccd1 _16615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ hold5663/X _13767_/A _13826_/X vssd1 vssd1 vccd1 vccd1 _13827_/Y sky130_fd_sc_hd__a21oi_1
X_17595_ _17721_/CLK _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16546_ _18198_/CLK _16546_/D vssd1 vssd1 vccd1 vccd1 _16546_/Q sky130_fd_sc_hd__dfxtp_1
X_13758_ _13779_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ hold2119/X hold3696/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16477_ _18362_/CLK _16477_/D vssd1 vssd1 vccd1 vccd1 _16477_/Q sky130_fd_sc_hd__dfxtp_1
X_13689_ _13791_/A _13689_/B vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _18216_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15428_ hold371/X _09367_/A _15479_/B1 _17346_/Q vssd1 vssd1 vccd1 vccd1 _15428_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18147_ _18153_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
X_15359_ hold460/X _15485_/A2 _15488_/A2 hold672/X _15358_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5907 hold6049/X vssd1 vssd1 vccd1 vccd1 _09447_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5918 _17540_/Q vssd1 vssd1 vccd1 vccd1 hold5918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5929 _17536_/Q vssd1 vssd1 vccd1 vccd1 hold5929/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 hold95/X vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold226 hold49/X vssd1 vssd1 vccd1 vccd1 input18/A sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _18078_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold237 hold731/X vssd1 vssd1 vccd1 vccd1 hold732/A sky130_fd_sc_hd__buf_4
X_09920_ hold3201/X hold4473/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__mux2_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _17875_/CLK _17029_/D vssd1 vssd1 vccd1 vccd1 _17029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout706 _07787_/Y vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09851_ _18352_/Q _16441_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__mux2_1
Xfanout717 _13037_/A vssd1 vssd1 vccd1 vccd1 _12444_/A sky130_fd_sc_hd__clkbuf_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout728 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15234_/C1 sky130_fd_sc_hd__buf_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _15473_/A vssd1 vssd1 vccd1 vccd1 _15186_/C1 sky130_fd_sc_hd__buf_4
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _12444_/A hold505/X vssd1 vssd1 vccd1 vccd1 _16020_/D sky130_fd_sc_hd__and2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09782_ hold3193/X _16418_/Q _10580_/C vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__mux2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08733_ hold312/X hold854/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold855/A sky130_fd_sc_hd__mux2_1
XFILLER_0_213_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08730_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _08685_/S sky130_fd_sc_hd__or2_2
XFILLER_0_178_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _15324_/A hold583/X vssd1 vssd1 vccd1 vccd1 _15921_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _15545_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09147_ hold2603/X _09164_/B _09146_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09078_ _15519_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ _15543_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_202_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 hold771/A vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold782 hold782/A vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _11136_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11040_/X sky130_fd_sc_hd__or2_1
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2150 _08036_/X vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 _14197_/X vssd1 vssd1 vccd1 vccd1 _17899_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 _18148_/Q vssd1 vssd1 vccd1 vccd1 hold2172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _07840_/X vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ hold2502/X hold3254/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_216_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _15825_/Q vssd1 vssd1 vccd1 vccd1 hold2194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1460 _18301_/Q vssd1 vssd1 vccd1 vccd1 hold1460/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14730_ _15231_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14730_/X sky130_fd_sc_hd__or2_1
Xhold1471 _15226_/X vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ hold1363/X _17138_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__mux2_1
Xhold1482 _15198_/X vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 _18391_/Q vssd1 vssd1 vccd1 vccd1 hold1493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ hold2407/X _14664_/B _14660_/Y _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14661_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ hold590/X hold4729/X _13793_/S vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _18377_/CLK _16400_/D vssd1 vssd1 vccd1 vccd1 _16400_/Q sky130_fd_sc_hd__dfxtp_1
X_13612_ hold4149/X _13802_/B _13611_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13612_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _11694_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14592_ _15201_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__or2_1
X_17380_ _17510_/CLK _17380_/D vssd1 vssd1 vccd1 vccd1 _17380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16331_ _18370_/CLK _16331_/D vssd1 vssd1 vccd1 vccd1 _16331_/Q sky130_fd_sc_hd__dfxtp_1
X_13543_ hold5703/X _13829_/B _13542_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13543_/X
+ sky130_fd_sc_hd__o211a_1
X_10755_ _11637_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _17496_/CLK _16262_/D vssd1 vssd1 vccd1 vccd1 _16262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ hold4413/X _13847_/B _13473_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10686_ _11643_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _15213_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__or2_1
X_18001_ _18064_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ hold607/X hold860/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold861/A sky130_fd_sc_hd__mux2_1
XFILLER_0_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16193_ _17478_/CLK _16193_/D vssd1 vssd1 vccd1 vccd1 _16193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15144_ hold1733/X _15167_/B _15143_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _17276_/Q _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _12234_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or2_1
X_15075_ _15183_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ hold1436/X hold3821/X _12302_/C vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14026_ _15533_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_457_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11238_ _12204_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ hold3604/X _11070_/A _11168_/X vssd1 vssd1 vccd1 vccd1 _11169_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _18410_/CLK _15977_/D vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _17748_/CLK _17716_/D vssd1 vssd1 vccd1 vccd1 _17716_/Q sky130_fd_sc_hd__dfxtp_1
X_14928_ _15197_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17647_ _17647_/CLK _17647_/D vssd1 vssd1 vccd1 vccd1 _17647_/Q sky130_fd_sc_hd__dfxtp_1
X_14859_ hold1791/X _14882_/B _14858_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14859_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_216_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _14328_/A hold2020/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_202_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17578_ _17703_/CLK _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ _18113_/CLK _16529_/D vssd1 vssd1 vccd1 vccd1 _16529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09001_ _12430_/A hold555/X vssd1 vssd1 vccd1 vccd1 _16117_/D sky130_fd_sc_hd__and2_1
XFILLER_0_6_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5704 _13543_/X vssd1 vssd1 vccd1 vccd1 _17634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5715 _17729_/Q vssd1 vssd1 vccd1 vccd1 hold5715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5726 _13507_/X vssd1 vssd1 vccd1 vccd1 _17622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5737 _17646_/Q vssd1 vssd1 vccd1 vccd1 hold5737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5748 _13537_/X vssd1 vssd1 vccd1 vccd1 _17632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5759 _17726_/Q vssd1 vssd1 vccd1 vccd1 hold5759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_198_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18380_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09903_ _11064_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout503 _10400_/S vssd1 vssd1 vccd1 vccd1 _10628_/C sky130_fd_sc_hd__clkbuf_8
Xfanout514 _10400_/S vssd1 vssd1 vccd1 vccd1 _10589_/C sky130_fd_sc_hd__clkbuf_8
Xfanout525 _09273_/S vssd1 vssd1 vccd1 vccd1 _09283_/S sky130_fd_sc_hd__buf_6
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout536 _08868_/X vssd1 vssd1 vccd1 vccd1 _12507_/A3 sky130_fd_sc_hd__buf_6
X_09834_ _09984_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_127_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17304_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout547 hold205/X vssd1 vssd1 vccd1 vccd1 _08390_/S sky130_fd_sc_hd__clkbuf_8
Xfanout558 hold239/X vssd1 vssd1 vccd1 vccd1 _08152_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout569 _07884_/Y vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__buf_8
XFILLER_0_225_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09765_ _09963_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08716_ _12404_/A hold880/X vssd1 vssd1 vccd1 vccd1 _15979_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09696_ _09984_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__or2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ hold578/X hold636/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ hold263/X hold318/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__mux2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10540_ hold4845/X _11180_/B _10539_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ hold4099/X _10571_/B _10470_/X _14827_/C1 vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _12213_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ _13190_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__or2_1
X_12141_ _13773_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12072_ _13773_/A _12072_/B vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__or2_1
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15900_ _17303_/CLK _15900_/D vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__dfxtp_1
X_11023_ hold5439/X _11198_/B _11022_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11023_/X
+ sky130_fd_sc_hd__o211a_1
X_16880_ _18049_/CLK _16880_/D vssd1 vssd1 vccd1 vccd1 _16880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _17722_/CLK _15831_/D vssd1 vssd1 vccd1 vccd1 _15831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _17501_/Q _12973_/X _12974_/S vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__mux2_1
X_15762_ _17681_/CLK _15762_/D vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 _08499_/X vssd1 vssd1 vccd1 vccd1 _15878_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ _18043_/CLK _17501_/D vssd1 vssd1 vccd1 vccd1 _17501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ hold3043/X _14714_/B _14712_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14713_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _13797_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__or2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _17199_/CLK _15693_/D vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _18456_/CLK _17432_/D vssd1 vssd1 vccd1 vccd1 _17432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_47_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_47_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14644_ _14984_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__or2_1
X_11856_ _13461_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ hold5142/X _11216_/B _10806_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__o211a_1
X_14575_ hold1865/X _14610_/B _14574_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14575_/X
+ sky130_fd_sc_hd__o211a_1
X_17363_ _17365_/CLK _17363_/D vssd1 vssd1 vccd1 vccd1 _17363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ hold4895/X _12234_/A _11786_/X vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16314_ _16323_/CLK _16314_/D vssd1 vssd1 vccd1 vccd1 _16314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10738_ hold5192/X _11216_/B _10737_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10738_/X
+ sky130_fd_sc_hd__o211a_1
X_13526_ hold2523/X hold3848/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17294_ _18410_/CLK _17294_/D vssd1 vssd1 vccd1 vccd1 hold670/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13457_ _15843_/Q _17606_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13458_/B sky130_fd_sc_hd__mux2_1
X_16245_ _17425_/CLK hold106/X vssd1 vssd1 vccd1 vccd1 _16245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10669_ hold3476/X _10019_/B _10668_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _10669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12408_ _12408_/A hold509/X vssd1 vssd1 vccd1 vccd1 _17297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ hold1735/X hold3629/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__mux2_1
X_16176_ _17482_/CLK _16176_/D vssd1 vssd1 vccd1 vccd1 _16176_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput106 hold5898/X vssd1 vssd1 vccd1 vccd1 ki sky130_fd_sc_hd__buf_12
XFILLER_0_140_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput117 hold5879/X vssd1 vssd1 vccd1 vccd1 hold5880/A sky130_fd_sc_hd__buf_6
XFILLER_0_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15127_ _15128_/A hold393/X vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__nor2_2
Xoutput128 hold5856/X vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_12
X_12339_ hold4952/X _12243_/A _12338_/X vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__a21oi_1
Xoutput139 _09339_/A vssd1 vssd1 vccd1 vccd1 load_data sky130_fd_sc_hd__buf_12
XFILLER_0_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3609 _17510_/Q vssd1 vssd1 vccd1 vccd1 hold3609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15058_ _15058_/A hold395/X vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_291_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2908 _14175_/X vssd1 vssd1 vccd1 vccd1 _17888_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2919 _18035_/Q vssd1 vssd1 vccd1 vccd1 hold2919/X sky130_fd_sc_hd__dlygate4sd3_1
X_14009_ hold2697/X _14038_/B _14008_/X _08131_/A vssd1 vssd1 vccd1 vccd1 _14009_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_220_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18113_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07880_ hold1436/X _07865_/B _07879_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _07880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ hold4809/X _10049_/B _09549_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09550_/X
+ sky130_fd_sc_hd__o211a_1
X_08501_ hold1744/X _08488_/B _08500_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _08501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09481_ _09482_/B _09484_/B _09481_/C vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ hold1929/X _08433_/B _08431_/Y _08391_/A vssd1 vssd1 vccd1 vccd1 _08432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08363_ _12657_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _15813_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ hold2038/X _08336_/A2 _08293_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _08294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_379_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17731_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5501 _17018_/Q vssd1 vssd1 vccd1 vccd1 hold5501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5512 _12244_/X vssd1 vssd1 vccd1 vccd1 _17238_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5523 _16818_/Q vssd1 vssd1 vccd1 vccd1 hold5523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5534 _11677_/X vssd1 vssd1 vccd1 vccd1 _17049_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4800 _10186_/X vssd1 vssd1 vccd1 vccd1 _16552_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5545 _17044_/Q vssd1 vssd1 vccd1 vccd1 hold5545/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_308_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17935_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4811 _16667_/Q vssd1 vssd1 vccd1 vccd1 hold4811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5556 _11278_/X vssd1 vssd1 vccd1 vccd1 _16916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4822 _09952_/X vssd1 vssd1 vccd1 vccd1 _16474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5567 _17076_/Q vssd1 vssd1 vccd1 vccd1 hold5567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4833 _16505_/Q vssd1 vssd1 vccd1 vccd1 hold4833/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5578 _11659_/X vssd1 vssd1 vccd1 vccd1 _17043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4844 _09664_/X vssd1 vssd1 vccd1 vccd1 _16378_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5589 _16750_/Q vssd1 vssd1 vccd1 vccd1 hold5589/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4855 _16381_/Q vssd1 vssd1 vccd1 vccd1 hold4855/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4866 _10171_/X vssd1 vssd1 vccd1 vccd1 _16547_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout300 _09987_/A vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__buf_4
Xhold4877 _16451_/Q vssd1 vssd1 vccd1 vccd1 hold4877/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout311 _10467_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__buf_4
XFILLER_0_160_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4888 _10714_/X vssd1 vssd1 vccd1 vccd1 _16728_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout322 _10470_/A vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__buf_4
Xhold4899 _16602_/Q vssd1 vssd1 vccd1 vccd1 hold4899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout333 fanout334/X vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__buf_4
Xfanout344 _09006_/S vssd1 vssd1 vccd1 vccd1 _09056_/S sky130_fd_sc_hd__buf_8
XFILLER_0_195_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout355 _08592_/S vssd1 vssd1 vccd1 vccd1 _08594_/S sky130_fd_sc_hd__buf_8
Xfanout366 hold734/X vssd1 vssd1 vccd1 vccd1 _15125_/B sky130_fd_sc_hd__buf_6
X_09817_ hold3802/X _10007_/B _09816_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09817_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout377 _14892_/B vssd1 vssd1 vccd1 vccd1 _14894_/B sky130_fd_sc_hd__buf_6
Xfanout388 _14680_/Y vssd1 vssd1 vccd1 vccd1 _14714_/B sky130_fd_sc_hd__buf_6
Xfanout399 _14446_/A2 vssd1 vssd1 vccd1 vccd1 _14433_/B sky130_fd_sc_hd__buf_6
XFILLER_0_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ hold5076/X _10034_/B _09747_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09748_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ hold3613/X _10577_/B _09678_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_95_wb_clk_i clkbuf_6_19_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18404_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ hold5002/X _12317_/B _11709_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12768_/A _12690_/B vssd1 vssd1 vccd1 vccd1 _17406_/D sky130_fd_sc_hd__and2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17469_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11641_ hold5158/X _11738_/B _11640_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _11641_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ _14360_/A _14360_/B vssd1 vssd1 vccd1 vccd1 _17977_/D sky130_fd_sc_hd__and2_1
XFILLER_0_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11572_ hold5557/X _11762_/B _11571_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13311_/A1 _13309_/X _13310_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13311_/X
+ sky130_fd_sc_hd__o211a_1
Xinput19 input19/A vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_10523_ hold1710/X _16665_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14291_ hold1753/X hold756/X _14290_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14291_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16030_ _17286_/CLK _16030_/D vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13242_ _17581_/Q _17115_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10454_ hold1843/X _16642_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _13172_/X hold3545/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10385_ hold1990/X hold3716/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ hold5356/X _13862_/B _12123_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12124_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17981_ _18459_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
X_12055_ hold4435/X _12365_/B _12054_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _12055_/X
+ sky130_fd_sc_hd__o211a_1
X_16932_ _18426_/CLK _16932_/D vssd1 vssd1 vccd1 vccd1 _16932_/Q sky130_fd_sc_hd__dfxtp_1
X_11006_ hold1682/X _16826_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__mux2_1
X_16863_ _18064_/CLK _16863_/D vssd1 vssd1 vccd1 vccd1 _16863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _17722_/CLK _15814_/D vssd1 vssd1 vccd1 vccd1 _15814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16794_ _18030_/CLK _16794_/D vssd1 vssd1 vccd1 vccd1 _16794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15745_ _17748_/CLK _15745_/D vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _12990_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _17495_/D sky130_fd_sc_hd__and2_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ hold5146/X _13798_/A2 _11907_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11908_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15676_ _17718_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12975_/A _12888_/B vssd1 vssd1 vccd1 vccd1 _17472_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17429_/CLK _17415_/D vssd1 vssd1 vccd1 vccd1 _17415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14627_ _14627_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14676_/B sky130_fd_sc_hd__or2_4
XFILLER_0_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18395_ _18395_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ hold5358/X _12314_/B _11838_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _17346_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 _17346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ hold690/X _14573_/B hold1218/X vssd1 vssd1 vccd1 vccd1 _14558_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _13713_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17277_ _17711_/CLK _17277_/D vssd1 vssd1 vccd1 vccd1 _17277_/Q sky130_fd_sc_hd__dfxtp_1
X_14489_ _15169_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14489_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16228_ _18456_/CLK _16228_/D vssd1 vssd1 vccd1 vccd1 _16228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4107 _17725_/Q vssd1 vssd1 vccd1 vccd1 hold4107/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_401_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17855_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4118 _15481_/X vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16159_ _17505_/CLK _16159_/D vssd1 vssd1 vccd1 vccd1 _16159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4129 _17659_/Q vssd1 vssd1 vccd1 vccd1 hold4129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3406 _09625_/X vssd1 vssd1 vccd1 vccd1 _16365_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08981_ hold263/X hold296/X _08993_/S vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__mux2_1
Xhold3417 _17595_/Q vssd1 vssd1 vccd1 vccd1 hold3417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3428 _17691_/Q vssd1 vssd1 vccd1 vccd1 hold3428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3439 _11140_/X vssd1 vssd1 vccd1 vccd1 _16870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2705 _18013_/Q vssd1 vssd1 vccd1 vccd1 hold2705/X sky130_fd_sc_hd__dlygate4sd3_1
X_07932_ _15555_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__or2_1
Xhold2716 _08400_/X vssd1 vssd1 vccd1 vccd1 _15830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2727 _15791_/Q vssd1 vssd1 vccd1 vccd1 hold2727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2738 _14195_/X vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 _09211_/X vssd1 vssd1 vccd1 vccd1 _16217_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ _14946_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09602_ hold1678/X hold3968/X _10004_/C vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07794_ _11158_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ _18246_/Q _13150_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _09463_/A _09461_/X _09484_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08415_ _15529_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ _15394_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _16284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ _14116_/A hold2611/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08277_ hold2564/X _08268_/B _08276_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08277_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6010 hold6034/X vssd1 vssd1 vccd1 vccd1 hold6010/X sky130_fd_sc_hd__buf_1
XFILLER_0_225_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6021 la_data_in[2] vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6032 _16316_/Q vssd1 vssd1 vccd1 vccd1 hold6032/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6043 la_data_in[13] vssd1 vssd1 vccd1 vccd1 hold6043/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5320 _16955_/Q vssd1 vssd1 vccd1 vccd1 hold5320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5331 _10333_/X vssd1 vssd1 vccd1 vccd1 _16601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_142_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18396_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5342 _17028_/Q vssd1 vssd1 vccd1 vccd1 hold5342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5353 _11362_/X vssd1 vssd1 vccd1 vccd1 _16944_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5364 _17212_/Q vssd1 vssd1 vccd1 vccd1 hold5364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4630 _16532_/Q vssd1 vssd1 vccd1 vccd1 hold4630/X sky130_fd_sc_hd__clkbuf_2
Xhold5375 _17198_/Q vssd1 vssd1 vccd1 vccd1 hold5375/X sky130_fd_sc_hd__dlygate4sd3_1
X_10170_ _10554_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__or2_1
Xhold4641 _17095_/Q vssd1 vssd1 vccd1 vccd1 hold4641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5386 _11305_/X vssd1 vssd1 vccd1 vccd1 _16925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4652 _10017_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5397 _17133_/Q vssd1 vssd1 vccd1 vccd1 hold5397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4663 _11781_/Y vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4674 _16909_/Q vssd1 vssd1 vccd1 vccd1 hold4674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3940 _17073_/Q vssd1 vssd1 vccd1 vccd1 hold3940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4685 _16342_/Q vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3951 _10327_/X vssd1 vssd1 vccd1 vccd1 _16599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4696 _12330_/Y vssd1 vssd1 vccd1 vccd1 _12331_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3962 _16576_/Q vssd1 vssd1 vccd1 vccd1 hold3962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3973 _10315_/X vssd1 vssd1 vccd1 vccd1 _16595_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3984 hold5869/X vssd1 vssd1 vccd1 vccd1 hold5870/A sky130_fd_sc_hd__buf_4
Xfanout152 _12827_/S vssd1 vssd1 vccd1 vccd1 _12914_/S sky130_fd_sc_hd__buf_6
Xfanout163 _12293_/B vssd1 vssd1 vccd1 vccd1 _13798_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3995 _12154_/X vssd1 vssd1 vccd1 vccd1 _17208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout174 _11150_/B vssd1 vssd1 vccd1 vccd1 _11617_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_227_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout185 _13777_/A2 vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout196 _12338_/B vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__buf_4
XFILLER_0_236_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13860_ hold3649/X _13788_/A _13859_/X vssd1 vssd1 vccd1 vccd1 _13860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12811_ hold2882/X hold3181/X _12913_/S vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13791_ _13791_/A _13791_/B vssd1 vssd1 vccd1 vccd1 _13791_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15530_ hold2959/X _15547_/B _15529_/X _12654_/A vssd1 vssd1 vccd1 vccd1 _15530_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _16245_/Q hold3195/X _12748_/S vssd1 vssd1 vccd1 vccd1 _12742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ hold723/X _09362_/D _09392_/D hold860/X _15460_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/D sky130_fd_sc_hd__a221o_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ hold2134/X hold3334/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17200_ _17200_/CLK _17200_/D vssd1 vssd1 vccd1 vccd1 _17200_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ hold1483/X hold5216/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__mux2_1
X_14412_ hold3112/X _14446_/A2 _14411_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14412_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18180_ _18180_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15392_ _15480_/A _15392_/B _15392_/C _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/X
+ sky130_fd_sc_hd__or4_1
X_17131_ _17195_/CLK _17131_/D vssd1 vssd1 vccd1 vccd1 _17131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14343_ hold915/X hold1397/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11555_ hold1620/X hold4493/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_231_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _10542_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or2_1
X_14274_ _15169_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
X_17062_ _17908_/CLK _17062_/D vssd1 vssd1 vccd1 vccd1 _17062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ hold1359/X _16986_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__and2_1
X_16013_ _18418_/CLK _16013_/D vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _10533_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ hold3604/X _13155_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ _10470_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__or2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ hold2403/X hold5156/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13199_/A1 _13085_/X _13086_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__o211a_1
X_17964_ _18050_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10533_/A _10299_/B vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12038_ hold2355/X hold4160/X _12362_/C vssd1 vssd1 vccd1 vccd1 _12039_/B sky130_fd_sc_hd__mux2_1
X_16915_ _17858_/CLK _16915_/D vssd1 vssd1 vccd1 vccd1 _16915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17895_ _17895_/CLK _17895_/D vssd1 vssd1 vccd1 vccd1 _17895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16846_ _18337_/CLK _16846_/D vssd1 vssd1 vccd1 vccd1 _16846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16777_ _18010_/CLK _16777_/D vssd1 vssd1 vccd1 vccd1 _16777_/Q sky130_fd_sc_hd__dfxtp_1
X_13989_ hold2104/X _13986_/B _13988_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _13989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15728_ _17667_/CLK _15728_/D vssd1 vssd1 vccd1 vccd1 _15728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _18447_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
X_15659_ _17171_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08200_ hold2638/X _08209_/B _08199_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08200_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09180_ _15509_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18378_ _18378_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__and2_1
X_17329_ _17329_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 _17329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08062_ _15521_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3203 _16499_/Q vssd1 vssd1 vccd1 vccd1 hold3203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3214 _14522_/X vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3225 _17474_/Q vssd1 vssd1 vccd1 vccd1 hold3225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3236 _18082_/Q vssd1 vssd1 vccd1 vccd1 hold3236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3247 _09996_/Y vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2502 _16171_/Q vssd1 vssd1 vccd1 vccd1 hold2502/X sky130_fd_sc_hd__dlygate4sd3_1
X_08964_ _09053_/A hold166/X vssd1 vssd1 vccd1 vccd1 _16099_/D sky130_fd_sc_hd__and2_1
Xhold3258 _12542_/X vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2513 _14275_/X vssd1 vssd1 vccd1 vccd1 _17936_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 _18176_/Q vssd1 vssd1 vccd1 vccd1 hold2524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 _17488_/Q vssd1 vssd1 vccd1 vccd1 hold3269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2535 _17517_/Q vssd1 vssd1 vccd1 vccd1 hold2535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1801 _18210_/Q vssd1 vssd1 vccd1 vccd1 hold1801/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2546 _18218_/Q vssd1 vssd1 vccd1 vccd1 hold2546/X sky130_fd_sc_hd__dlygate4sd3_1
X_07915_ hold2667/X _07918_/B _07914_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07915_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1812 _15184_/X vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08895_ _15324_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _16065_/D sky130_fd_sc_hd__and2_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2557 _15727_/Q vssd1 vssd1 vccd1 vccd1 hold2557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _18033_/Q vssd1 vssd1 vccd1 vccd1 hold1823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 _16152_/Q vssd1 vssd1 vccd1 vccd1 hold2568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _09439_/X vssd1 vssd1 vccd1 vccd1 _16305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 _16220_/Q vssd1 vssd1 vccd1 vccd1 hold2579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1845 _17945_/Q vssd1 vssd1 vccd1 vccd1 hold1845/X sky130_fd_sc_hd__dlygate4sd3_1
X_07846_ hold1350/X _07869_/B _07845_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _07846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1856 _14633_/X vssd1 vssd1 vccd1 vccd1 _18107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _18346_/Q vssd1 vssd1 vccd1 vccd1 hold1867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 _09336_/X vssd1 vssd1 vccd1 vccd1 _16278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 la_data_in[8] vssd1 vssd1 vccd1 vccd1 hold1889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ _09918_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ _09447_/A _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09456_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_394_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17804_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09378_ hold458/X _09367_/A _09386_/D hold651/X vssd1 vssd1 vccd1 vccd1 _09378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _15553_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_323_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17777_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_152_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _11631_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _11658_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11271_/X sky130_fd_sc_hd__or2_1
X_13010_ hold1404/X _13003_/Y _13009_/X _12531_/A vssd1 vssd1 vccd1 vccd1 _13010_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5150 _17228_/Q vssd1 vssd1 vccd1 vccd1 hold5150/X sky130_fd_sc_hd__dlygate4sd3_1
X_10222_ hold4909/X _10649_/B _10221_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5161 _11905_/X vssd1 vssd1 vccd1 vccd1 _17125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5172 _17623_/Q vssd1 vssd1 vccd1 vccd1 hold5172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5183 _10378_/X vssd1 vssd1 vccd1 vccd1 _16616_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5194 _16590_/Q vssd1 vssd1 vccd1 vccd1 hold5194/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4460 _11020_/X vssd1 vssd1 vccd1 vccd1 _16830_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10153_ hold4921/X _10631_/B _10152_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10153_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4471 _16963_/Q vssd1 vssd1 vccd1 vccd1 hold4471/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4482 _09634_/X vssd1 vssd1 vccd1 vccd1 _16368_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4493 _17009_/Q vssd1 vssd1 vccd1 vccd1 hold4493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3770 _17399_/Q vssd1 vssd1 vccd1 vccd1 hold3770/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14961_ hold1857/X _14952_/B _14960_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14961_/X
+ sky130_fd_sc_hd__o211a_1
X_10084_ hold5693/X _10598_/B _10083_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _10084_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3781 _17413_/Q vssd1 vssd1 vccd1 vccd1 hold3781/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3792 _13872_/Y vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_4
XFILLER_0_227_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16700_ _18212_/CLK _16700_/D vssd1 vssd1 vccd1 vccd1 _16700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13912_ _14862_/A hold2155/X hold124/X vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__mux2_1
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ _17680_/CLK _17680_/D vssd1 vssd1 vccd1 vccd1 _17680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _15231_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16631_ _16631_/CLK _16631_/D vssd1 vssd1 vccd1 vccd1 _16631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13843_ _13873_/A _13843_/B vssd1 vssd1 vccd1 vccd1 _17734_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _18208_/CLK _16562_/D vssd1 vssd1 vccd1 vccd1 _16562_/Q sky130_fd_sc_hd__dfxtp_1
X_10986_ _11082_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10986_/X sky130_fd_sc_hd__or2_1
X_13774_ hold4093/X _13868_/B _13773_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _13774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18301_ _18309_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15513_ _15513_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__or2_1
X_12725_ hold3676/X _12724_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__mux2_1
X_16493_ _18396_/CLK _16493_/D vssd1 vssd1 vccd1 vccd1 _16493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18232_ _18232_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
X_15444_ _15482_/A _15444_/B vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__and2_1
X_12656_ hold3661/X _12655_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18163_ _18163_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _12057_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ hold422/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__or2_1
X_12587_ hold3300/X _12586_/X _12965_/S vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _17178_/CLK _17114_/D vssd1 vssd1 vccd1 vccd1 _17114_/Q sky130_fd_sc_hd__dfxtp_1
X_14326_ _14774_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18094_ _18222_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11538_ _11637_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold408 hold408/A vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold419 hold419/A vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17045_ _17901_/CLK _17045_/D vssd1 vssd1 vccd1 vccd1 _17045_/Q sky130_fd_sc_hd__dfxtp_1
X_14257_ hold2496/X _14266_/B _14256_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14257_/X
+ sky130_fd_sc_hd__o211a_1
X_11469_ _11667_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _13201_/X _13207_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17544_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14188_ _15207_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _13138_/X _16910_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_238_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17947_ _18429_/CLK hold757/X vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1108 hold1108/A vssd1 vssd1 vccd1 vccd1 hold1108/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 _17780_/Q vssd1 vssd1 vccd1 vccd1 hold1119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _12418_/A hold882/X vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17878_ _17878_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_6_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16829_ _18030_/CLK _16829_/D vssd1 vssd1 vccd1 vccd1 _16829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09301_ _15523_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ hold331/X hold533/X vssd1 vssd1 vccd1 vccd1 hold534/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09163_ hold2626/X _09164_/B _09162_/Y _12912_/A vssd1 vssd1 vccd1 vccd1 _09163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ _15519_/A hold1040/X hold240/X vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09094_ _15535_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ _14894_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold920 hold955/X vssd1 vssd1 vccd1 vccd1 hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold931 hold931/A vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold942 hold947/X vssd1 vssd1 vccd1 vccd1 hold948/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 hold964/A vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3000 _18205_/Q vssd1 vssd1 vccd1 vccd1 hold3000/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3011 _14426_/X vssd1 vssd1 vccd1 vccd1 _18009_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3022 _07848_/X vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 _18345_/Q vssd1 vssd1 vccd1 vccd1 hold3033/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 input48/X vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__buf_1
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _13102_/A _09918_/A _09995_/X vssd1 vssd1 vccd1 vccd1 _09996_/Y sky130_fd_sc_hd__a21oi_1
Xhold3044 _14713_/X vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3055 _18117_/Q vssd1 vssd1 vccd1 vccd1 hold3055/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2310 _15570_/Q vssd1 vssd1 vccd1 vccd1 hold2310/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3066 _09097_/X vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 _15655_/Q vssd1 vssd1 vccd1 vccd1 hold2321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3077 hold5826/X vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2332 _13961_/X vssd1 vssd1 vccd1 vccd1 _17785_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08947_ hold47/X hold846/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__mux2_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3088 _18056_/Q vssd1 vssd1 vccd1 vccd1 hold3088/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2343 _15596_/Q vssd1 vssd1 vccd1 vccd1 hold2343/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2354 _14783_/X vssd1 vssd1 vccd1 vccd1 _18180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3099 _17976_/Q vssd1 vssd1 vccd1 vccd1 hold3099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 _18151_/Q vssd1 vssd1 vccd1 vccd1 hold2365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 _17855_/Q vssd1 vssd1 vccd1 vccd1 hold1620/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2376 _08249_/X vssd1 vssd1 vccd1 vccd1 _15759_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 _08465_/X vssd1 vssd1 vccd1 vccd1 _15861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 _18147_/Q vssd1 vssd1 vccd1 vccd1 hold1642/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2387 _17939_/Q vssd1 vssd1 vccd1 vccd1 hold2387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2398 _14587_/X vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ hold88/X _16057_/Q _08932_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1653 _08422_/X vssd1 vssd1 vccd1 vccd1 _15841_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1664 _18132_/Q vssd1 vssd1 vccd1 vccd1 hold1664/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1675 _08235_/X vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1686 _16252_/Q vssd1 vssd1 vccd1 vccd1 hold1686/X sky130_fd_sc_hd__dlygate4sd3_1
X_07829_ _14843_/A hold202/X vssd1 vssd1 vccd1 vccd1 _07829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_224_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 _18001_/Q vssd1 vssd1 vccd1 vccd1 hold1697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ hold5615/X _11768_/B _10839_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _10840_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ hold3515/X _10019_/B _10770_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12510_ _14556_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12510_/Y sky130_fd_sc_hd__nor2_1
X_13490_ hold1379/X _17617_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12441_ hold498/X hold771/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold772/A sky130_fd_sc_hd__mux2_1
XFILLER_0_192_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15160_ hold1573/X _15167_/B _15159_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _15160_/X
+ sky130_fd_sc_hd__o211a_1
X_12372_ hold3736/X _13782_/A _12371_/X vssd1 vssd1 vccd1 vccd1 _12372_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11323_ hold4471/X _11801_/B _11322_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11323_/X
+ sky130_fd_sc_hd__o211a_1
X_14111_ hold1759/X _14148_/B _14110_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14111_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15091_ _15199_/A hold734/X vssd1 vssd1 vccd1 vccd1 _15091_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14042_ _14328_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__or2_1
X_11254_ hold5395/X _11732_/B _11253_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10205_ hold3097/X hold4936/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11185_ _11218_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _16885_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4290 _12187_/X vssd1 vssd1 vccd1 vccd1 _17219_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17801_ _17821_/CLK _17801_/D vssd1 vssd1 vccd1 vccd1 _17801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10136_ hold1797/X _16536_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__mux2_1
XTAP_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ _18415_/CLK _15993_/D vssd1 vssd1 vccd1 vccd1 hold611/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _17732_/CLK _17732_/D vssd1 vssd1 vccd1 vccd1 _17732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ _16513_/Q _10565_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10067_/X sky130_fd_sc_hd__and3_1
X_14944_ _15213_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ _17695_/CLK _17663_/D vssd1 vssd1 vccd1 vccd1 _17663_/Q sky130_fd_sc_hd__dfxtp_1
X_14875_ hold1914/X _14882_/B _14874_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16614_ _18170_/CLK _16614_/D vssd1 vssd1 vccd1 vccd1 _16614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _17729_/Q _13832_/B _13826_/C vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__and3_1
X_17594_ _17722_/CLK _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_245_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18144_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _18230_/CLK _16545_/D vssd1 vssd1 vccd1 vccd1 _16545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ hold2436/X _17706_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__mux2_1
X_10969_ hold5066/X _11159_/B _10968_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _10969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12708_ _12768_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _17412_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16476_ _18387_/CLK _16476_/D vssd1 vssd1 vccd1 vccd1 _16476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ hold1742/X hold4372/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ _18215_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ hold660/X _09392_/B _09392_/C hold217/X vssd1 vssd1 vccd1 vccd1 _15427_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _12810_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _17389_/D sky130_fd_sc_hd__and2_1
XFILLER_0_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _18178_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15358_ hold547/X _15484_/A2 _09392_/D hold574/X vssd1 vssd1 vccd1 vccd1 _15358_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5908 hold6041/X vssd1 vssd1 vccd1 vccd1 _09463_/C sky130_fd_sc_hd__buf_1
XFILLER_0_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__buf_2
Xhold5919 _16915_/Q vssd1 vssd1 vccd1 vccd1 hold5919/X sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ hold2921/X hold756/X _14308_/X _14442_/C1 vssd1 vssd1 vccd1 vccd1 _14309_/X
+ sky130_fd_sc_hd__o211a_1
X_18077_ _18202_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ hold404/X _15485_/A2 _15488_/A2 hold370/X _15288_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold227 input18/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__buf_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__clkbuf_4
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _17897_/CLK _17028_/D vssd1 vssd1 vccd1 vccd1 _17028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 _15374_/A vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__clkbuf_4
X_09850_ hold5176/X _11177_/B _09849_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09850_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 _13037_/A vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__clkbuf_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout729 _14915_/C1 vssd1 vssd1 vccd1 vccd1 _15052_/A sky130_fd_sc_hd__buf_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ hold215/X hold504/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ hold3657/X _10049_/B _09780_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09781_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _09055_/A hold794/X vssd1 vssd1 vccd1 vccd1 _15986_/D sky130_fd_sc_hd__and2_1
XFILLER_0_217_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ _13043_/C hold990/X vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_1
XFILLER_0_240_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08594_ hold150/X hold582/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold583/A sky130_fd_sc_hd__mux2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09215_ hold2027/X _09216_/B _09214_/Y _12894_/A vssd1 vssd1 vccd1 vccd1 _09215_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09146_ _15529_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_228_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09077_ hold2049/X _09119_/A2 _09076_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18039_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08028_ hold2321/X _08029_/B _08027_/Y _08137_/A vssd1 vssd1 vccd1 vccd1 _08028_/X
+ sky130_fd_sc_hd__o211a_1
Xhold750 hold750/A vssd1 vssd1 vccd1 vccd1 input55/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 la_data_in[28] vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold783 hold783/A vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold794 hold794/A vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ hold4737/X _10601_/B _09978_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09979_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 next_key vssd1 vssd1 vccd1 vccd1 hold2140/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2151 _15871_/Q vssd1 vssd1 vccd1 vccd1 hold2151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2162 _15591_/Q vssd1 vssd1 vccd1 vccd1 hold2162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2173 _14717_/X vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12990_/A _12990_/B vssd1 vssd1 vccd1 vccd1 _17506_/D sky130_fd_sc_hd__and2_1
XFILLER_0_207_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2184 _16168_/Q vssd1 vssd1 vccd1 vccd1 hold2184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1450 _18053_/Q vssd1 vssd1 vccd1 vccd1 hold1450/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2195 _15863_/Q vssd1 vssd1 vccd1 vccd1 hold2195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _15035_/X vssd1 vssd1 vccd1 vccd1 _15036_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ hold5114/X _12347_/B _11940_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _11941_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1472 _17883_/Q vssd1 vssd1 vccd1 vccd1 hold1472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 _17878_/Q vssd1 vssd1 vccd1 vccd1 hold1483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _15222_/X vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14660_ _14946_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__nand2_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ hold3436/X _12347_/B _11871_/X _08125_/A vssd1 vssd1 vccd1 vccd1 _11872_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_37_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_37_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13611_ _13713_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ hold1307/X hold4509/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__mux2_1
X_14591_ hold2280/X _14610_/B _14590_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16330_ _18273_/CLK _16330_/D vssd1 vssd1 vccd1 vccd1 _16330_/Q sky130_fd_sc_hd__dfxtp_1
X_13542_ _13734_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ hold1753/X hold4211/X _11729_/C vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _17365_/CLK _16261_/D vssd1 vssd1 vccd1 vccd1 _16261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13473_ _13746_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__or2_1
X_10685_ hold2113/X hold3591/X _11738_/C vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__mux2_1
X_18000_ _18059_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ hold1851/X _15219_/B _15211_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15212_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12424_ _12424_/A hold655/X vssd1 vssd1 vccd1 vccd1 _17305_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16192_ _17878_/CLK _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _15197_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _13825_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _17275_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _17772_/Q hold4895/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__mux2_1
X_15074_ hold733/X hold393/X vssd1 vssd1 vccd1 vccd1 hold734/A sky130_fd_sc_hd__or2_1
X_12286_ hold4964/X _12317_/B _12285_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _12286_/X
+ sky130_fd_sc_hd__o211a_1
X_11237_ hold1972/X hold4683/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__mux2_1
X_14025_ hold2414/X _14040_/B _14024_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _14025_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11168_ _16880_/Q _11168_/B _11168_/C vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__and3_1
XTAP_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10563_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _17298_/CLK _15976_/D vssd1 vssd1 vccd1 vccd1 hold899/A sky130_fd_sc_hd__dfxtp_1
X_11099_ hold2886/X hold4861/X _11192_/C vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_234_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _17747_/CLK _17715_/D vssd1 vssd1 vccd1 vccd1 _17715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14927_ hold1070/X _14946_/B _14926_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_426_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17199_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17646_ _17731_/CLK _17646_/D vssd1 vssd1 vccd1 vccd1 _17646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _15197_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13809_ _17563_/Q _13713_/A _13808_/X vssd1 vssd1 vccd1 vccd1 _13809_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17577_ _17641_/CLK _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
X_14789_ _14789_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14830_/B sky130_fd_sc_hd__or2_4
X_16528_ _18208_/CLK _16528_/D vssd1 vssd1 vccd1 vccd1 _16528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ _18364_/CLK _16459_/D vssd1 vssd1 vccd1 vccd1 _16459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09000_ hold554/X _16117_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold555/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18129_ _18181_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5705 _17730_/Q vssd1 vssd1 vccd1 vccd1 hold5705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5716 _13732_/X vssd1 vssd1 vccd1 vccd1 _17697_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5727 _17699_/Q vssd1 vssd1 vccd1 vccd1 hold5727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5738 _13483_/X vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5749 _17741_/Q vssd1 vssd1 vccd1 vccd1 hold5749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09902_ hold2766/X hold5110/X _11159_/C vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__mux2_1
Xfanout504 _10400_/S vssd1 vssd1 vccd1 vccd1 _10997_/S sky130_fd_sc_hd__clkbuf_8
Xfanout515 _10613_/C vssd1 vssd1 vccd1 vccd1 _10619_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 hold534/X vssd1 vssd1 vccd1 vccd1 _09273_/S sky130_fd_sc_hd__clkbuf_8
X_09833_ hold1867/X hold3386/X _10007_/C vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__mux2_1
Xfanout537 _08868_/X vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_226_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout548 _08299_/B vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__buf_8
Xfanout559 _08100_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__buf_6
XFILLER_0_158_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ hold3151/X _16412_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08715_ hold222/X hold879/X _08727_/S vssd1 vssd1 vccd1 vccd1 hold880/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_167_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18395_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09695_ hold2507/X _16389_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _12438_/A hold406/X vssd1 vssd1 vccd1 vccd1 _15945_/D sky130_fd_sc_hd__and2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08577_ _15364_/A hold696/X vssd1 vssd1 vccd1 vccd1 _15912_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ _10470_/A _10470_/B vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ hold1227/X _09177_/A2 _09128_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ hold1256/X _17204_/Q _13868_/C vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_241_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12071_ hold2042/X hold3434/X _12251_/S vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 hold591/A vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _11103_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _17721_/CLK _15830_/D vssd1 vssd1 vccd1 vccd1 _15830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_239_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _17680_/CLK _15761_/D vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfxtp_1
X_12973_ _16165_/Q _17502_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux2_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1280 _14883_/X vssd1 vssd1 vccd1 vccd1 _18228_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _18043_/CLK _17500_/D vssd1 vssd1 vccd1 vccd1 _17500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14712_ _15105_/A _14730_/B vssd1 vssd1 vccd1 vccd1 _14712_/X sky130_fd_sc_hd__or2_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 _17774_/Q vssd1 vssd1 vccd1 vccd1 hold1291/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ hold1132/X hold5024/X _13412_/S vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _17260_/CLK _15692_/D vssd1 vssd1 vccd1 vccd1 _15692_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17431_/CLK _17431_/D vssd1 vssd1 vccd1 vccd1 _17431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ hold1771/X _14666_/B _14642_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14643_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ hold2572/X hold3627/X _13556_/S vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__mux2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10806_ _11121_/A _10806_/B vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__or2_1
X_17362_ _17510_/CLK _17362_/D vssd1 vssd1 vccd1 vccd1 _17362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14574_ _14968_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _17086_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _16323_/CLK _16313_/D vssd1 vssd1 vccd1 vccd1 _16313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13525_ hold4073/X _13802_/B _13524_/X _13714_/C1 vssd1 vssd1 vccd1 vccd1 _13525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17293_ _17293_/CLK _17293_/D vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__dfxtp_1
X_10737_ _11121_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _17425_/CLK hold448/X vssd1 vssd1 vccd1 vccd1 _16244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13456_ hold4321/X _13856_/B _13455_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _11136_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ hold454/X hold508/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold509/A sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _18460_/CLK _16175_/D vssd1 vssd1 vccd1 vccd1 _16175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ hold3545/X _10563_/A _10598_/X vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__a21oi_1
X_13387_ hold5757/X _13817_/B _13386_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _13387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput107 hold4271/X vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ hold3033/X _15113_/B _15125_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15126_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput118 hold5854/X vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_12
Xoutput129 hold5851/X vssd1 vssd1 vccd1 vccd1 hold5852/A sky130_fd_sc_hd__buf_6
X_12338_ _17270_/Q _12338_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15057_ hold181/X _18312_/Q _15071_/S vssd1 vssd1 vccd1 vccd1 hold395/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ hold2890/X _17247_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2909 _18061_/Q vssd1 vssd1 vccd1 vccd1 hold2909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14008_ _14116_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_260_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15959_ _17321_/CLK _15959_/D vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08500_ _14894_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ hold850/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__and2_1
XFILLER_0_231_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ _15004_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__nand2_1
X_17629_ _17722_/CLK _17629_/D vssd1 vssd1 vccd1 vccd1 _17629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08362_ _15531_/A hold2290/X hold134/X vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08293_ _14403_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5502 _11488_/X vssd1 vssd1 vccd1 vccd1 _16986_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5513 _17012_/Q vssd1 vssd1 vccd1 vccd1 hold5513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5524 _10888_/X vssd1 vssd1 vccd1 vccd1 _16786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5535 _16747_/Q vssd1 vssd1 vccd1 vccd1 hold5535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4801 _16474_/Q vssd1 vssd1 vccd1 vccd1 hold4801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5546 _11566_/X vssd1 vssd1 vccd1 vccd1 _17012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4812 _10435_/X vssd1 vssd1 vccd1 vccd1 _16635_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5557 _17046_/Q vssd1 vssd1 vccd1 vccd1 hold5557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4823 _16792_/Q vssd1 vssd1 vccd1 vccd1 hold4823/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5568 _11662_/X vssd1 vssd1 vccd1 vccd1 _17044_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4834 _09949_/X vssd1 vssd1 vccd1 vccd1 _16473_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5579 _16876_/Q vssd1 vssd1 vccd1 vccd1 hold5579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4845 _16702_/Q vssd1 vssd1 vccd1 vccd1 hold4845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4856 _09577_/X vssd1 vssd1 vccd1 vccd1 _16349_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4867 _16700_/Q vssd1 vssd1 vccd1 vccd1 hold4867/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout301 _09843_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_4
Xhold4878 _09787_/X vssd1 vssd1 vccd1 vccd1 _16419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout312 _11097_/A vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__buf_2
XFILLER_0_160_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout323 _09564_/A vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4889 _16628_/Q vssd1 vssd1 vccd1 vccd1 hold4889/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout334 _09493_/Y vssd1 vssd1 vccd1 vccd1 fanout334/X sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_348_wb_clk_i clkbuf_6_42_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17641_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout345 _08997_/S vssd1 vssd1 vccd1 vccd1 _08993_/S sky130_fd_sc_hd__buf_8
XFILLER_0_195_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout356 _08536_/S vssd1 vssd1 vccd1 vccd1 _08592_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09816_ _09936_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__or2_1
Xfanout367 hold765/X vssd1 vssd1 vccd1 vccd1 _15113_/B sky130_fd_sc_hd__buf_8
Xfanout378 _14842_/Y vssd1 vssd1 vccd1 vccd1 _14882_/B sky130_fd_sc_hd__buf_8
Xfanout389 _14676_/B vssd1 vssd1 vccd1 vccd1 _14678_/B sky130_fd_sc_hd__buf_6
XFILLER_0_94_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09747_ _09843_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09678_ _10488_/A _09678_/B vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08629_ hold346/X hold588/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__mux2_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11643_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _11667_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11571_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13310_ _13310_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_64_wb_clk_i clkbuf_6_24_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18012_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10522_ _10616_/A _11198_/B _10521_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14290_ _15185_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13241_ _13241_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__and2_1
XFILLER_0_165_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10453_ hold3958/X _10646_/B _10452_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10384_ hold4847/X _11177_/B _10383_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10384_/X
+ sky130_fd_sc_hd__o211a_1
X_13172_ hold3691/X _13171_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ _12261_/A _12123_/B vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_241_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17980_ _18012_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12054_ _12246_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__or2_1
X_16931_ _17777_/CLK _16931_/D vssd1 vssd1 vccd1 vccd1 _16931_/Q sky130_fd_sc_hd__dfxtp_1
X_11005_ hold4861/X _11180_/B _11004_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _11005_/X
+ sky130_fd_sc_hd__o211a_1
X_16862_ _17999_/CLK _16862_/D vssd1 vssd1 vccd1 vccd1 _16862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15813_ _18448_/CLK _15813_/D vssd1 vssd1 vccd1 vccd1 _15813_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout890 hold525/X vssd1 vssd1 vccd1 vccd1 _14854_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_232_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16793_ _17994_/CLK _16793_/D vssd1 vssd1 vccd1 vccd1 _16793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15744_ _17683_/CLK _15744_/D vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ hold3244/X _12955_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12956_/X sky130_fd_sc_hd__mux2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11907_ _13797_/A _11907_/B vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__or2_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15675_ _17898_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12887_ hold3301/X _12886_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12888_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_200_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17429_/CLK _17414_/D vssd1 vssd1 vccd1 vccd1 _17414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14626_ _14627_/A hold393/X vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nor2_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _18394_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11838_ _12219_/A _11838_/B vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__or2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17345_ _17346_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _17345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ hold690/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_173_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ hold5004/X _11694_/A _11768_/X vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13508_ hold2037/X _17623_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17276_ _17276_/CLK _17276_/D vssd1 vssd1 vccd1 vccd1 _17276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14488_ hold2620/X _14487_/B _14487_/Y _14356_/A vssd1 vssd1 vccd1 vccd1 _14488_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16227_ _17459_/CLK _16227_/D vssd1 vssd1 vccd1 vccd1 _16227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ hold2327/X hold5743/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13440_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _17505_/CLK hold969/X vssd1 vssd1 vccd1 vccd1 hold968/A sky130_fd_sc_hd__dfxtp_1
Xhold4108 hold5895/X vssd1 vssd1 vccd1 vccd1 hold5896/A sky130_fd_sc_hd__buf_6
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4119 _16836_/Q vssd1 vssd1 vccd1 vccd1 hold4119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _15217_/A _15113_/B vssd1 vssd1 vccd1 vccd1 _15109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3407 _17456_/Q vssd1 vssd1 vccd1 vccd1 hold3407/X sky130_fd_sc_hd__dlygate4sd3_1
X_08980_ _13037_/A hold657/X vssd1 vssd1 vccd1 vccd1 _16107_/D sky130_fd_sc_hd__and2_1
XFILLER_0_224_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16089_ _16089_/CLK _16089_/D vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3418 _13330_/X vssd1 vssd1 vccd1 vccd1 _17563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3429 _13618_/X vssd1 vssd1 vccd1 vccd1 _17659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2706 _14434_/X vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_441_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17658_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07931_ hold2816/X _07924_/B _07930_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _07931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2717 _15635_/Q vssd1 vssd1 vccd1 vccd1 hold2717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 _08316_/X vssd1 vssd1 vccd1 vccd1 _15791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2739 _16191_/Q vssd1 vssd1 vccd1 vccd1 hold2739/X sky130_fd_sc_hd__dlygate4sd3_1
X_07862_ hold2669/X _07865_/B _07861_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07862_/X
+ sky130_fd_sc_hd__o211a_1
X_09601_ hold3408/X _10025_/B _09600_/X _15454_/A vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ hold5913/X _07788_/A hold1412/X _14556_/A vssd1 vssd1 vccd1 vccd1 _07793_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09532_ hold3960/X _10010_/B _09531_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09463_ _09463_/A _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09472_/D
+ sky130_fd_sc_hd__and4_2
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ hold2327/X _08433_/B _08413_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08414_/X
+ sky130_fd_sc_hd__o211a_1
X_09394_ hold5884/A _15481_/B1 _09393_/X _15490_/A1 vssd1 vssd1 vccd1 vccd1 _09394_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _08389_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _15804_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08276_ _15555_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6000 _16149_/Q vssd1 vssd1 vccd1 vccd1 hold6000/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6011 data_in[7] vssd1 vssd1 vccd1 vccd1 hold593/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6022 la_data_in[24] vssd1 vssd1 vccd1 vccd1 hold716/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6033 data_in[28] vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6044 data_in[4] vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5310 _16878_/Q vssd1 vssd1 vccd1 vccd1 hold5310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5321 _11299_/X vssd1 vssd1 vccd1 vccd1 _16923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5332 _17094_/Q vssd1 vssd1 vccd1 vccd1 hold5332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5343 _11518_/X vssd1 vssd1 vccd1 vccd1 _16996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5354 _16585_/Q vssd1 vssd1 vccd1 vccd1 hold5354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4620 _10635_/Y vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5365 _12070_/X vssd1 vssd1 vccd1 vccd1 _17180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4631 _10605_/Y vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5376 _12028_/X vssd1 vssd1 vccd1 vccd1 _17166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4642 _12294_/Y vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5387 _16394_/Q vssd1 vssd1 vccd1 vccd1 hold5387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5398 _11833_/X vssd1 vssd1 vccd1 vccd1 _17101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4653 _17102_/Q vssd1 vssd1 vccd1 vccd1 hold4653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4664 _16723_/Q vssd1 vssd1 vccd1 vccd1 hold4664/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3930 _16996_/Q vssd1 vssd1 vccd1 vccd1 hold3930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4675 _11736_/Y vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4686 _10035_/Y vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_182_wb_clk_i clkbuf_6_51_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3941 _11653_/X vssd1 vssd1 vccd1 vccd1 _17041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3952 _16705_/Q vssd1 vssd1 vccd1 vccd1 hold3952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4697 _16910_/Q vssd1 vssd1 vccd1 vccd1 hold4697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3963 _10162_/X vssd1 vssd1 vccd1 vccd1 _16544_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_111_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3974 _16879_/Q vssd1 vssd1 vccd1 vccd1 hold3974/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout153 _12974_/S vssd1 vssd1 vccd1 vccd1 _12827_/S sky130_fd_sc_hd__buf_4
Xhold3985 _15363_/X vssd1 vssd1 vccd1 vccd1 _15364_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout164 _13808_/B vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__buf_4
Xhold3996 _17034_/Q vssd1 vssd1 vccd1 vccd1 hold3996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout175 _11150_/B vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout186 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _13777_/A2 sky130_fd_sc_hd__buf_4
Xfanout197 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _12338_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12810_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _17446_/D sky130_fd_sc_hd__and2_1
XFILLER_0_236_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13790_ hold2761/X hold4330/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13791_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_232_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _17423_/D sky130_fd_sc_hd__and2_1
XFILLER_0_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _07805_/A _15477_/A2 _09392_/A hold836/X vssd1 vssd1 vccd1 vccd1 _15460_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12672_ _12810_/A _12672_/B vssd1 vssd1 vccd1 vccd1 _17400_/D sky130_fd_sc_hd__and2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14984_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__or2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ hold5012/X _12299_/B _11622_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _11623_/X
+ sky130_fd_sc_hd__o211a_1
X_15391_ _16303_/Q _09362_/A _09392_/B hold846/X _15390_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_154_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _17161_/CLK _17130_/D vssd1 vssd1 vccd1 vccd1 _17130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ _14388_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _17968_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ hold5423/X _11732_/B _11553_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10505_ hold1298/X hold4061/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__mux2_1
X_17061_ _17907_/CLK _17061_/D vssd1 vssd1 vccd1 vccd1 _17061_/Q sky130_fd_sc_hd__dfxtp_1
X_14273_ hold2432/X _14272_/B _14272_/Y _13917_/A vssd1 vssd1 vccd1 vccd1 _14273_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ hold5525/X _12338_/B _11484_/X _14131_/C1 vssd1 vssd1 vccd1 vccd1 _11485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _18418_/CLK _16012_/D vssd1 vssd1 vccd1 vccd1 _16012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ _13217_/X _13223_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17546_/D sky130_fd_sc_hd__o21a_1
X_10436_ hold2770/X hold3954/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ _13154_/X _16912_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_237_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ hold3084/X _16613_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ hold4927/X _13811_/B _12105_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _12106_/X
+ sky130_fd_sc_hd__o211a_1
X_13086_ _13086_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__or2_1
X_10298_ hold3043/X hold5194/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10299_/B sky130_fd_sc_hd__mux2_1
X_17963_ _17994_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12037_ hold3464/X _13871_/B _12036_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12037_/X
+ sky130_fd_sc_hd__o211a_1
X_16914_ _17889_/CLK _16914_/D vssd1 vssd1 vccd1 vccd1 _16914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17894_ _17894_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _18046_/CLK _16845_/D vssd1 vssd1 vccd1 vccd1 _16845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16776_ _18041_/CLK _16776_/D vssd1 vssd1 vccd1 vccd1 _16776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _14328_/A _13996_/B vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _17730_/CLK _15727_/D vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfxtp_1
X_12939_ _12999_/A _12939_/B vssd1 vssd1 vccd1 vccd1 _17489_/D sky130_fd_sc_hd__and2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_238_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18446_ _18448_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
X_15658_ _17170_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ hold2252/X _14612_/B _14608_/Y _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14609_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18377_ _18377_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15589_ _17274_/CLK _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08130_ _14529_/A hold1609/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__mux2_1
X_17328_ _17344_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _17328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ hold1314/X _08097_/A2 _08060_/X _15500_/A vssd1 vssd1 vccd1 vccd1 _08061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _18428_/CLK _17259_/D vssd1 vssd1 vccd1 vccd1 _17259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3204 _09931_/X vssd1 vssd1 vccd1 vccd1 _16467_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3215 _17502_/Q vssd1 vssd1 vccd1 vccd1 hold3215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3226 _12893_/X vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3237 _14581_/X vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08963_ hold118/X hold165/X _08963_/S vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3248 _16328_/Q vssd1 vssd1 vccd1 vccd1 _13094_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2503 _09113_/X vssd1 vssd1 vccd1 vccd1 _16171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3259 _17351_/Q vssd1 vssd1 vccd1 vccd1 hold3259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _17894_/Q vssd1 vssd1 vccd1 vccd1 hold2514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2525 _14775_/X vssd1 vssd1 vccd1 vccd1 _18176_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2536 _13018_/X vssd1 vssd1 vccd1 vccd1 _17517_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07914_ _15537_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07914_/X sky130_fd_sc_hd__or2_1
Xhold1802 _14847_/X vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2547 _14863_/X vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1813 _18105_/Q vssd1 vssd1 vccd1 vccd1 hold1813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ hold271/X hold396/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2558 _08182_/X vssd1 vssd1 vccd1 vccd1 _15727_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 _14476_/X vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 _09075_/X vssd1 vssd1 vccd1 vccd1 _16152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1835 _18370_/Q vssd1 vssd1 vccd1 vccd1 hold1835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1846 _14295_/X vssd1 vssd1 vccd1 vccd1 _17945_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07845_ _14517_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07845_/X sky130_fd_sc_hd__or2_1
Xhold1857 _18265_/Q vssd1 vssd1 vccd1 vccd1 hold1857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 _15130_/X vssd1 vssd1 vccd1 vccd1 _18346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1879 _18048_/Q vssd1 vssd1 vccd1 vccd1 hold1879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09515_ _18240_/Q _13102_/A _10019_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09444_/X _09446_/B _09484_/B vssd1 vssd1 vccd1 vccd1 _16308_/D sky130_fd_sc_hd__and3b_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09377_ hold5858/A _09342_/B _09342_/Y _09376_/X _12412_/A vssd1 vssd1 vccd1 vccd1
+ _09377_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08328_ hold1395/X _08323_/B _08327_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08259_ hold1742/X _08263_/A2 _08258_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_363_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17711_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11270_ hold1507/X hold4907/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5140 _16697_/Q vssd1 vssd1 vccd1 vccd1 hold5140/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ _10533_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__or2_1
Xhold5151 _12118_/X vssd1 vssd1 vccd1 vccd1 _17196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5162 _16386_/Q vssd1 vssd1 vccd1 vccd1 hold5162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5173 _13414_/X vssd1 vssd1 vccd1 vccd1 _17591_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5184 _17062_/Q vssd1 vssd1 vccd1 vccd1 hold5184/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5195 _10204_/X vssd1 vssd1 vccd1 vccd1 _16558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4450 _13393_/X vssd1 vssd1 vccd1 vccd1 _17584_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ _10536_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or2_1
Xhold4461 _17747_/Q vssd1 vssd1 vccd1 vccd1 hold4461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4472 _11323_/X vssd1 vssd1 vccd1 vccd1 _16931_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4483 _17618_/Q vssd1 vssd1 vccd1 vccd1 hold4483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4494 _11461_/X vssd1 vssd1 vccd1 vccd1 _16977_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3760 _17409_/Q vssd1 vssd1 vccd1 vccd1 hold3760/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _15121_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__or2_1
X_10083_ _10191_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10083_/X sky130_fd_sc_hd__or2_1
Xhold3771 _12668_/X vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3782 _16441_/Q vssd1 vssd1 vccd1 vccd1 hold3782/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3793 _16629_/Q vssd1 vssd1 vccd1 vccd1 hold3793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _13911_/A _13911_/B vssd1 vssd1 vccd1 vccd1 _17761_/D sky130_fd_sc_hd__and2_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ hold1214/X _14882_/B _14890_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14891_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ _18198_/CLK _16630_/D vssd1 vssd1 vccd1 vccd1 _16630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ hold3702/X _13746_/A _13841_/X vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16561_ _18181_/CLK _16561_/D vssd1 vssd1 vccd1 vccd1 _16561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13773_ _13773_/A _13773_/B vssd1 vssd1 vccd1 vccd1 _13773_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ hold1693/X _16819_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18300_ _18300_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ hold1261/X _15507_/Y _15511_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _15512_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ hold2205/X hold3508/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16492_ _18303_/CLK _16492_/D vssd1 vssd1 vccd1 vccd1 _16492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18231_ _18231_/CLK _18231_/D vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15481_/A1 _15435_/X _15442_/X _15481_/B1 hold5882/A vssd1 vssd1 vccd1 vccd1
+ _15443_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12655_ hold2844/X hold3466/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18162_ _18182_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ hold1557/X hold4491/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__mux2_1
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12586_ hold2033/X hold3275/X _12601_/S vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17113_ _17113_/CLK _17113_/D vssd1 vssd1 vccd1 vccd1 _17113_/Q sky130_fd_sc_hd__dfxtp_1
X_14325_ hold1988/X _14326_/B _14324_/Y _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14325_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18093_ _18213_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
X_11537_ hold2858/X hold4179/X _11729_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17044_ _17858_/CLK _17044_/D vssd1 vssd1 vccd1 vccd1 _17044_/Q sky130_fd_sc_hd__dfxtp_1
X_14256_ _14758_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__or2_1
X_11468_ hold1549/X hold5497/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _13311_/A1 _13205_/X _13206_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13207_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _10497_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14187_ hold2514/X _14202_/B _14186_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11399_ hold1287/X hold5385/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _17568_/Q _17102_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13138_/X sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13068_/X hold4795/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17946_ _18012_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _08354_/X vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17877_ _17877_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16828_ _18061_/CLK _16828_/D vssd1 vssd1 vccd1 vccd1 _16828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_232_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16759_ _18124_/CLK _16759_/D vssd1 vssd1 vccd1 vccd1 _16759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ hold2622/X _09338_/A2 _09299_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ hold1881/X _09216_/B _09230_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _09231_/X
+ sky130_fd_sc_hd__o211a_1
X_18429_ _18429_/CLK hold693/X vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09162_ _15545_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08113_ _13927_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09093_ hold2991/X _09106_/B _09092_/X _12969_/A vssd1 vssd1 vccd1 vccd1 _09093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ hold1410/X _08033_/B _08043_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _08044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 hold910/A vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold921 hold956/X vssd1 vssd1 vccd1 vccd1 hold957/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_222_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold943 hold949/X vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__buf_2
Xhold3001 _14835_/X vssd1 vssd1 vccd1 vccd1 _18205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/A vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 hold976/A vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3012 _17856_/Q vssd1 vssd1 vccd1 vccd1 hold3012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 hold998/A vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__buf_8
Xhold3023 _18439_/Q vssd1 vssd1 vccd1 vccd1 hold3023/X sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _16489_/Q _10013_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__and3_1
Xhold3034 _15126_/X vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3045 _16268_/Q vssd1 vssd1 vccd1 vccd1 hold3045/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2300 _15782_/Q vssd1 vssd1 vccd1 vccd1 hold2300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3056 _14653_/X vssd1 vssd1 vccd1 vccd1 _18117_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2311 _07850_/X vssd1 vssd1 vccd1 vccd1 _15570_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2322 _08028_/X vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08946_ _12426_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _16090_/D sky130_fd_sc_hd__and2_1
Xhold3067 _18140_/Q vssd1 vssd1 vccd1 vccd1 hold3067/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3078 _13047_/X vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2333 _15730_/Q vssd1 vssd1 vccd1 vccd1 hold2333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3089 _14524_/X vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2344 _07905_/X vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 _15658_/Q vssd1 vssd1 vccd1 vccd1 hold2355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 _17870_/Q vssd1 vssd1 vccd1 vccd1 hold1610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 _14723_/X vssd1 vssd1 vccd1 vccd1 _18151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1621 _14105_/X vssd1 vssd1 vccd1 vccd1 _17855_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1632 _17923_/Q vssd1 vssd1 vccd1 vccd1 hold1632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08877_ _15364_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _16056_/D sky130_fd_sc_hd__and2_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2377 _16195_/Q vssd1 vssd1 vccd1 vccd1 hold2377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 _14715_/X vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 _14281_/X vssd1 vssd1 vccd1 vccd1 _17939_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2399 _15603_/Q vssd1 vssd1 vccd1 vccd1 hold2399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1654 _17904_/Q vssd1 vssd1 vccd1 vccd1 hold1654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1665 _14685_/X vssd1 vssd1 vccd1 vccd1 _18132_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1676 _18100_/Q vssd1 vssd1 vccd1 vccd1 hold1676/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _14556_/A hold531/A _14555_/C vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__or3_1
XFILLER_0_93_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 _15864_/Q vssd1 vssd1 vccd1 vccd1 hold1687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_27_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_27_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold1698 _14410_/X vssd1 vssd1 vccd1 vccd1 _18001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _11136_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09429_ _07804_/A _09472_/A _15344_/A _09428_/X vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ _12444_/A hold599/X vssd1 vssd1 vccd1 vccd1 _17313_/D sky130_fd_sc_hd__and2_1
XFILLER_0_125_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ _17281_/Q _13877_/B _13877_/C vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14110_ _14164_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _11706_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__or2_1
X_15090_ hold1646/X _15113_/B _15089_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ hold2529/X _14040_/B _14040_/Y _13909_/A vssd1 vssd1 vccd1 vccd1 _14041_/X
+ sky130_fd_sc_hd__o211a_1
X_11253_ _11553_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10204_ hold5194/X _10625_/B _10203_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ hold4678/X _11121_/A _11183_/X vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__a21oi_1
XTAP_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4280 _10756_/X vssd1 vssd1 vccd1 vccd1 _16742_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17800_ _17860_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ hold3752/X _10637_/B _10134_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _10135_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4291 hold5845/X vssd1 vssd1 vccd1 vccd1 hold5846/A sky130_fd_sc_hd__buf_4
XTAP_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ _17334_/CLK _15992_/D vssd1 vssd1 vccd1 vccd1 hold722/A sky130_fd_sc_hd__dfxtp_1
XTAP_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3590 _13809_/Y vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14943_ hold1827/X _14946_/B _14942_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _14943_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10066_ _10603_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _16512_/D sky130_fd_sc_hd__nor2_1
X_17731_ _17731_/CLK _17731_/D vssd1 vssd1 vccd1 vccd1 _17731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14874_ _15213_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__or2_1
X_17662_ _17666_/CLK _17662_/D vssd1 vssd1 vccd1 vccd1 _17662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16613_ _18201_/CLK _16613_/D vssd1 vssd1 vccd1 vccd1 _16613_/Q sky130_fd_sc_hd__dfxtp_1
X_13825_ _13825_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _17728_/D sky130_fd_sc_hd__nor2_1
X_17593_ _17721_/CLK _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ _18228_/CLK _16544_/D vssd1 vssd1 vccd1 vccd1 _16544_/Q sky130_fd_sc_hd__dfxtp_1
X_13756_ hold4366/X _13880_/B _13755_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10968_ _11064_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _10968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12707_ hold3786/X _12706_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__mux2_1
X_16475_ _18322_/CLK _16475_/D vssd1 vssd1 vccd1 vccd1 _16475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ hold3490/X _13880_/B _13686_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13687_/X
+ sky130_fd_sc_hd__o211a_1
X_10899_ _11103_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15426_ _17318_/Q _09357_/A _09392_/A hold848/X vssd1 vssd1 vccd1 vccd1 _15426_/X
+ sky130_fd_sc_hd__a22o_1
X_18214_ _18214_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_285_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18287_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12638_ hold3331/X _12637_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15357_ hold424/X _15487_/A2 _15484_/B1 hold494/X _15356_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/B sky130_fd_sc_hd__a221o_1
X_18145_ _18209_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_214_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ hold3488/X _12568_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5909 hold6032/X vssd1 vssd1 vccd1 vccd1 _09472_/C sky130_fd_sc_hd__buf_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _15529_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__or2_1
X_18076_ _18202_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
X_15288_ hold491/X _15484_/A2 _09392_/D hold303/X vssd1 vssd1 vccd1 vccd1 _15288_/X
+ sky130_fd_sc_hd__a22o_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold50/X vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__buf_4
XFILLER_0_22_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17027_ _17905_/CLK _17027_/D vssd1 vssd1 vccd1 vccd1 _17027_/Q sky130_fd_sc_hd__dfxtp_1
X_14239_ hold1658/X _14266_/B _14238_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__buf_1
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 _15374_/A vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__buf_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 _07787_/Y vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_237_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _12444_/A hold585/X vssd1 vssd1 vccd1 vccd1 _16019_/D sky130_fd_sc_hd__and2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _10470_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ hold554/X hold793/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold794/A sky130_fd_sc_hd__mux2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _18026_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_1411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08662_ _12418_/A hold700/X vssd1 vssd1 vccd1 vccd1 _15953_/D sky130_fd_sc_hd__and2_1
XFILLER_0_205_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08593_ _12412_/A hold908/X vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _15543_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_174_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ hold975/X _09164_/B _09144_/X _12990_/A vssd1 vssd1 vccd1 vccd1 hold976/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ _15517_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08027_ _15541_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold740 hold740/A vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold751 input55/X vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold762 hold762/A vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 hold773/A vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold784 hold784/A vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/A vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17515_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _10488_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__or2_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2130 _15607_/Q vssd1 vssd1 vccd1 vccd1 hold2130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2141 hold2141/A vssd1 vssd1 vccd1 vccd1 input69/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08929_ _15304_/A hold833/X vssd1 vssd1 vccd1 vccd1 _16082_/D sky130_fd_sc_hd__and2_1
Xhold2152 _08485_/X vssd1 vssd1 vccd1 vccd1 _15871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2163 _07895_/X vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2174 _15834_/Q vssd1 vssd1 vccd1 vccd1 hold2174/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1440 input62/X vssd1 vssd1 vccd1 vccd1 hold1440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2185 _09107_/X vssd1 vssd1 vccd1 vccd1 _16168_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 _14518_/X vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2196 _08469_/X vssd1 vssd1 vccd1 vccd1 _15863_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ _12261_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__or2_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1462 _15789_/Q vssd1 vssd1 vccd1 vccd1 hold1462/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1473 _14165_/X vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1484 _14153_/X vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _15777_/Q vssd1 vssd1 vccd1 vccd1 hold1495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _12231_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__or2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ hold2896/X _17657_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ hold5541/X _11753_/B _10821_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _10822_/X
+ sky130_fd_sc_hd__o211a_1
X_14590_ _14984_/A _14602_/B vssd1 vssd1 vccd1 vccd1 _14590_/X sky130_fd_sc_hd__or2_1
XFILLER_0_200_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13541_ _15819_/Q _17634_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10753_ hold5481/X _11156_/B _10752_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _17496_/CLK _16260_/D vssd1 vssd1 vccd1 vccd1 _16260_/Q sky130_fd_sc_hd__dfxtp_1
X_13472_ hold2079/X hold3484/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__mux2_1
X_10684_ hold5589/X _11201_/B _10683_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15211_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15211_/X sky130_fd_sc_hd__or2_1
X_12423_ hold228/X hold654/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold655/A sky130_fd_sc_hd__mux2_1
XFILLER_0_180_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16191_ _17478_/CLK _16191_/D vssd1 vssd1 vccd1 vccd1 _16191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ hold5989/X _15165_/B hold1031/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15142_/X
+ sky130_fd_sc_hd__o211a_1
X_12354_ hold4729/X _13794_/A _12353_/X vssd1 vssd1 vccd1 vccd1 _12354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11305_ hold5385/X _12329_/B _11304_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15073_ hold733/X hold393/X vssd1 vssd1 vccd1 vccd1 hold765/A sky130_fd_sc_hd__nor2_1
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__or2_1
X_14024_ _15531_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14024_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ hold5122/X _12308_/B _11235_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11236_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _12310_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _16879_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ hold1956/X hold3545/X _10580_/C vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__mux2_1
XTAP_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _18408_/CLK _15975_/D vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__dfxtp_1
X_11098_ _11192_/A _11192_/B _11097_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _11098_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _17746_/CLK _17714_/D vssd1 vssd1 vccd1 vccd1 _17714_/Q sky130_fd_sc_hd__dfxtp_1
X_10049_ _16507_/Q _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__and3_1
X_14926_ _15195_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17645_ _17677_/CLK _17645_/D vssd1 vssd1 vccd1 vccd1 _17645_/Q sky130_fd_sc_hd__dfxtp_1
X_14857_ hold1298/X _14880_/B _14856_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _13808_/A _13808_/B _13808_/C vssd1 vssd1 vccd1 vccd1 _13808_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14788_ _14789_/A hold392/X vssd1 vssd1 vccd1 vccd1 _14788_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_133_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17576_ _17738_/CLK _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
X_16527_ _18159_/CLK _16527_/D vssd1 vssd1 vccd1 vccd1 _16527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13739_ hold1567/X _17700_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _18395_/CLK _16458_/D vssd1 vssd1 vccd1 vccd1 _16458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15409_ hold193/X _15485_/A2 _15488_/A2 hold615/X _15408_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16389_ _17534_/CLK _16389_/D vssd1 vssd1 vccd1 vccd1 _16389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18128_ _18180_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5706 _13735_/X vssd1 vssd1 vccd1 vccd1 _17698_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5717 _17697_/Q vssd1 vssd1 vccd1 vccd1 hold5717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5728 _13642_/X vssd1 vssd1 vccd1 vccd1 _17667_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5739 _17635_/Q vssd1 vssd1 vccd1 vccd1 hold5739/X sky130_fd_sc_hd__dlygate4sd3_1
X_18059_ _18059_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ hold3375/X _10013_/B _09900_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09901_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout505 _10400_/S vssd1 vssd1 vccd1 vccd1 _10640_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout516 _10613_/C vssd1 vssd1 vccd1 vccd1 _10637_/C sky130_fd_sc_hd__clkbuf_8
X_09832_ hold5597/X _09832_/A2 _09831_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _09832_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout527 _09220_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__buf_4
Xfanout538 _08858_/S vssd1 vssd1 vccd1 vccd1 _08866_/S sky130_fd_sc_hd__buf_8
XFILLER_0_226_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout549 _08336_/A2 vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__buf_6
X_09763_ hold3662/X _10565_/B _09762_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09763_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ _12408_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _15978_/D sky130_fd_sc_hd__and2_1
XFILLER_0_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09694_ hold4097/X _11159_/B _09693_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08645_ hold263/X hold405/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold406/A sky130_fd_sc_hd__mux2_1
XFILLER_0_96_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08576_ hold607/X hold695/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__mux2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_136_wb_clk_i clkbuf_6_29_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16148_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09128_ hold999/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09059_ _09063_/A hold295/X vssd1 vssd1 vccd1 vccd1 _16146_/D sky130_fd_sc_hd__and2_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ hold5364/X _13862_/B _12069_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12070_/X
+ sky130_fd_sc_hd__o211a_1
Xhold570 hold570/A vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold581 hold581/A vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold592 hold592/A vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ hold2917/X _16831_/Q _11198_/C vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _17647_/CLK _15760_/D vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12975_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _17500_/D sky130_fd_sc_hd__and2_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 _07887_/X vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14711_ hold3095/X _14714_/B _14710_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14711_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_213_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1281 _17953_/Q vssd1 vssd1 vccd1 vccd1 hold1281/X sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ hold5186/X _12308_/B _11922_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11923_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1292 _18452_/Q vssd1 vssd1 vccd1 vccd1 hold1292/X sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ _17260_/CLK _15691_/D vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _15197_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _18455_/CLK _17430_/D vssd1 vssd1 vccd1 vccd1 _17430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ hold4087/X _13868_/B _11853_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11854_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ hold1988/X hold5078/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__mux2_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ hold238/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14602_/B sky130_fd_sc_hd__nand2_4
X_17361_ _17510_/CLK _17361_/D vssd1 vssd1 vccd1 vccd1 _17361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11785_ _12340_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _17085_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16312_ _16312_/CLK _16312_/D vssd1 vssd1 vccd1 vccd1 _16312_/Q sky130_fd_sc_hd__dfxtp_1
X_13524_ _13713_/A _13524_/B vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__or2_1
X_17292_ _17327_/CLK _17292_/D vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__dfxtp_1
X_10736_ hold1720/X hold4707/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16243_ _17689_/CLK _16243_/D vssd1 vssd1 vccd1 vccd1 _16243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13455_ _13761_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ hold1769/X _16713_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12406_ _15324_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _17296_/D sky130_fd_sc_hd__and2_1
XFILLER_0_125_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16174_ _17496_/CLK _16174_/D vssd1 vssd1 vccd1 vccd1 _16174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13386_ _13767_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__or2_1
X_10598_ _16690_/Q _10598_/B _11096_/S vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _15233_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput108 hold5836/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_12
X_12337_ _13873_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _17269_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput119 hold5882/X vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_239_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15056_ _15056_/A hold742/X vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12268_ hold4121/X _13871_/B _12267_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _12268_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14007_ hold1783/X _14038_/B _14006_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _14007_/X
+ sky130_fd_sc_hd__o211a_1
X_11219_ _16897_/Q _11789_/B _11219_/C vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__and3_1
X_12199_ hold4994/X _12293_/B _12198_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _12199_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput90 _13265_/A vssd1 vssd1 vccd1 vccd1 output90/X sky130_fd_sc_hd__buf_6
XFILLER_0_207_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15958_ _17321_/CLK _15958_/D vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__dfxtp_1
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ _18240_/Q _14896_/Y hold526/X _15394_/A vssd1 vssd1 vccd1 vccd1 hold527/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15889_ _17334_/CLK _15889_/D vssd1 vssd1 vccd1 vccd1 hold630/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ hold2128/X _08433_/B _08429_/Y _13750_/C1 vssd1 vssd1 vccd1 vccd1 _08430_/X
+ sky130_fd_sc_hd__o211a_1
X_17628_ _17723_/CLK _17628_/D vssd1 vssd1 vccd1 vccd1 _17628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08361_ _12738_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _17719_/CLK _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08292_ hold2660/X _08336_/A2 _08291_/X _13483_/C1 vssd1 vssd1 vccd1 vccd1 _08292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5503 _16744_/Q vssd1 vssd1 vccd1 vccd1 hold5503/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5514 _11470_/X vssd1 vssd1 vccd1 vccd1 _16980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5525 _17017_/Q vssd1 vssd1 vccd1 vccd1 hold5525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5536 _10675_/X vssd1 vssd1 vccd1 vccd1 _16715_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4802 _09856_/X vssd1 vssd1 vccd1 vccd1 _16442_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5547 _17050_/Q vssd1 vssd1 vccd1 vccd1 hold5547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4813 _16692_/Q vssd1 vssd1 vccd1 vccd1 hold4813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5558 _11572_/X vssd1 vssd1 vccd1 vccd1 _17014_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4824 _10810_/X vssd1 vssd1 vccd1 vccd1 _16760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5569 _16952_/Q vssd1 vssd1 vccd1 vccd1 hold5569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4835 _16583_/Q vssd1 vssd1 vccd1 vccd1 hold4835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4846 _10540_/X vssd1 vssd1 vccd1 vccd1 _16670_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4857 _16925_/Q vssd1 vssd1 vccd1 vccd1 hold4857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4868 _10534_/X vssd1 vssd1 vccd1 vccd1 _16668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout302 _11061_/A vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__buf_4
Xhold4879 _16587_/Q vssd1 vssd1 vccd1 vccd1 hold4879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout313 fanout334/X vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout324 _09564_/A vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__buf_4
Xfanout335 _12508_/B vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__buf_4
XFILLER_0_201_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout346 _08963_/S vssd1 vssd1 vccd1 vccd1 _08997_/S sky130_fd_sc_hd__buf_8
X_09815_ hold2308/X _16429_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout357 _15521_/B vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__buf_4
XFILLER_0_201_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout368 hold765/X vssd1 vssd1 vccd1 vccd1 _15111_/B sky130_fd_sc_hd__clkbuf_8
Xfanout379 _14842_/Y vssd1 vssd1 vccd1 vccd1 _14880_/B sky130_fd_sc_hd__buf_6
XFILLER_0_199_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09746_ _18317_/Q hold3365/X _10034_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_388_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17170_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ hold1601/X _16383_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_317_wb_clk_i clkbuf_6_47_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18068_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ _09055_/A hold459/X vssd1 vssd1 vccd1 vccd1 _15936_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_234_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08559_ _12418_/A hold841/X vssd1 vssd1 vccd1 vccd1 _15903_/D sky130_fd_sc_hd__and2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11570_ hold2550/X hold5437/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _11103_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ _13233_/X _13239_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ _10998_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13171_ _13170_/X hold4907/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__mux2_1
X_10383_ _11082_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18043_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12122_ hold1371/X _17198_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12053_ hold1410/X _17175_/Q _12365_/C vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__mux2_1
X_16930_ _17808_/CLK _16930_/D vssd1 vssd1 vccd1 vccd1 _16930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _11100_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__or2_1
X_16861_ _18062_/CLK _16861_/D vssd1 vssd1 vccd1 vccd1 _16861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout880 hold1723/X vssd1 vssd1 vccd1 vccd1 hold1724/A sky130_fd_sc_hd__buf_6
XFILLER_0_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout891 hold926/X vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__buf_12
X_15812_ _17422_/CLK _15812_/D vssd1 vssd1 vccd1 vccd1 _15812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16792_ _18200_/CLK _16792_/D vssd1 vssd1 vccd1 vccd1 _16792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12955_ hold2797/X _17496_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__mux2_1
X_15743_ _17746_/CLK _15743_/D vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11906_ hold1098/X _17126_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__mux2_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _18462_/A vssd1 vssd1 vccd1 vccd1 _18462_/X sky130_fd_sc_hd__buf_1
XFILLER_0_59_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15674_ _17166_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12886_ hold1614/X hold3173/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__mux2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17413_ _17413_/CLK _17413_/D vssd1 vssd1 vccd1 vccd1 _17413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14625_ hold3047/X _14612_/B _14624_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14625_/X
+ sky130_fd_sc_hd__o211a_1
X_11837_ hold2106/X hold4691/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18393_ _18393_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17344_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _17344_/Q sky130_fd_sc_hd__dfxtp_1
X_14556_ _14556_/A hold531/A hold391/A vssd1 vssd1 vccd1 vccd1 hold392/A sky130_fd_sc_hd__or3_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11768_ _17080_/Q _11768_/B _11768_/C vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ _11103_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__or2_1
X_13507_ hold5725/X _13817_/B _13506_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13507_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14487_ _15547_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__nand2_1
X_17275_ _17741_/CLK _17275_/D vssd1 vssd1 vccd1 vccd1 _17275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ hold2218/X _17057_/Q _12365_/C vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13438_ hold5697/X _13829_/B _13437_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _13438_/X
+ sky130_fd_sc_hd__o211a_1
X_16226_ _18432_/CLK _16226_/D vssd1 vssd1 vccd1 vccd1 _16226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16157_ _17496_/CLK _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/Q sky130_fd_sc_hd__dfxtp_1
X_13369_ hold3529/X _13777_/A2 _13368_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13369_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4109 _15490_/X vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15108_ hold2234/X _15111_/B _15107_/Y _15186_/C1 vssd1 vssd1 vccd1 vccd1 _15108_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ _18410_/CLK _16088_/D vssd1 vssd1 vccd1 vccd1 hold518/A sky130_fd_sc_hd__dfxtp_1
Xhold3408 _16389_/Q vssd1 vssd1 vccd1 vccd1 hold3408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3419 _17459_/Q vssd1 vssd1 vccd1 vccd1 hold3419/X sky130_fd_sc_hd__dlygate4sd3_1
X_15039_ hold944/X hold1005/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__mux2_1
X_07930_ _15553_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2707 _17879_/Q vssd1 vssd1 vccd1 vccd1 hold2707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2718 _07985_/X vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2729 _15564_/Q vssd1 vssd1 vccd1 vccd1 hold2729/X sky130_fd_sc_hd__dlygate4sd3_1
X_07861_ _15539_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__or2_1
XFILLER_0_235_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09600_ _09984_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__or2_1
X_07792_ _18458_/Q vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _09933_/A _09531_/B vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_410_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17885_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09462_ _09461_/X _09484_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _16314_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_52_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08413_ _14862_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09393_ _07805_/Y _09362_/A _09369_/D _09392_/X vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_175_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08344_ _14794_/A hold1352/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ hold2650/X _08268_/B _08274_/X _13714_/C1 vssd1 vssd1 vccd1 vccd1 _08275_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6001 _18246_/Q vssd1 vssd1 vccd1 vccd1 hold6001/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6012 _18403_/Q vssd1 vssd1 vccd1 vccd1 hold6012/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6023 _16307_/Q vssd1 vssd1 vccd1 vccd1 hold6023/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6034 _18413_/Q vssd1 vssd1 vccd1 vccd1 hold6034/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6045 _16536_/Q vssd1 vssd1 vccd1 vccd1 hold6045/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5300 _16748_/Q vssd1 vssd1 vccd1 vccd1 hold5300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5311 _11068_/X vssd1 vssd1 vccd1 vccd1 _16846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5322 _16502_/Q vssd1 vssd1 vccd1 vccd1 hold5322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5333 _12292_/X vssd1 vssd1 vccd1 vccd1 _17254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5344 _16557_/Q vssd1 vssd1 vccd1 vccd1 hold5344/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4610 _16353_/Q vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5355 _10189_/X vssd1 vssd1 vccd1 vccd1 _16553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4621 _16539_/Q vssd1 vssd1 vccd1 vccd1 hold4621/X sky130_fd_sc_hd__buf_1
Xhold5366 _17168_/Q vssd1 vssd1 vccd1 vccd1 hold5366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4632 _16726_/Q vssd1 vssd1 vccd1 vccd1 hold4632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5377 _16973_/Q vssd1 vssd1 vccd1 vccd1 hold5377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5388 _09616_/X vssd1 vssd1 vccd1 vccd1 _16362_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4643 _17566_/Q vssd1 vssd1 vccd1 vccd1 hold4643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5399 _16396_/Q vssd1 vssd1 vccd1 vccd1 hold5399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4654 _12315_/Y vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3920 _16606_/Q vssd1 vssd1 vccd1 vccd1 hold3920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4665 _11178_/Y vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4676 _16730_/Q vssd1 vssd1 vccd1 vccd1 hold4676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3931 _11422_/X vssd1 vssd1 vccd1 vccd1 _16964_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4687 _16526_/Q vssd1 vssd1 vccd1 vccd1 hold4687/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3942 _17594_/Q vssd1 vssd1 vccd1 vccd1 hold3942/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3953 _10549_/X vssd1 vssd1 vccd1 vccd1 _16673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4698 _11739_/Y vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3964 _16326_/Q vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__buf_1
Xhold3975 _11071_/X vssd1 vssd1 vccd1 vccd1 _16847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout154 _12986_/S vssd1 vssd1 vccd1 vccd1 _12926_/S sky130_fd_sc_hd__buf_6
XFILLER_0_227_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3986 _16462_/Q vssd1 vssd1 vccd1 vccd1 hold3986/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout165 _13817_/B vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__buf_4
Xfanout176 _11150_/B vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__buf_4
Xhold3997 _11536_/X vssd1 vssd1 vccd1 vccd1 _17002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout187 _12347_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__buf_4
Xfanout198 _11210_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__buf_4
X_09729_ _11106_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_151_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18418_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ hold3199/X _12739_/X _12749_/S vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__mux2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ hold3795/X _12670_/X _12773_/S vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ hold1697/X _14446_/A2 _14409_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14410_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11712_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ hold759/X _09367_/A _09392_/A hold852/X vssd1 vssd1 vccd1 vccd1 _15390_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ _14968_/A hold1666/X hold333/X vssd1 vssd1 vccd1 vccd1 _14341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11553_ _11553_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ hold4869/X _11180_/B _10503_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o211a_1
X_17060_ _17908_/CLK _17060_/D vssd1 vssd1 vccd1 vccd1 _17060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14272_ _14774_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_150_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _12243_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16011_ _18300_/CLK _16011_/D vssd1 vssd1 vccd1 vccd1 hold385/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13223_ _13311_/A1 _13221_/X _13222_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ hold4811/X _10625_/B _10434_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ _17570_/Q _17104_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
X_10366_ hold3651/X _11180_/B _10365_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10366_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _13716_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13084_/X hold3543/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _17994_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
X_10297_ hold5312/X _10619_/B _10296_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10297_/X
+ sky130_fd_sc_hd__o211a_1
X_12036_ _12267_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__or2_1
X_16913_ _17855_/CLK _16913_/D vssd1 vssd1 vccd1 vccd1 _16913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_239_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18216_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17893_ _17970_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16844_ _18045_/CLK _16844_/D vssd1 vssd1 vccd1 vccd1 _16844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ _18010_/CLK _16775_/D vssd1 vssd1 vccd1 vccd1 _16775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ hold2494/X _13986_/B _13986_/Y _13921_/A vssd1 vssd1 vccd1 vccd1 _13987_/X
+ sky130_fd_sc_hd__o211a_1
X_15726_ _17695_/CLK _15726_/D vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ hold3267/X _12937_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12938_/X sky130_fd_sc_hd__mux2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18445_ _18445_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
X_15657_ _17266_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ hold3303/X _12868_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_186_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ _14878_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _18376_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15588_ _17236_/CLK _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ _17327_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _17327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539_ _15545_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _15519_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17258_ _17258_/CLK _17258_/D vssd1 vssd1 vccd1 vccd1 _17258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ _17446_/CLK _16209_/D vssd1 vssd1 vccd1 vccd1 _16209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17189_ _17189_/CLK _17189_/D vssd1 vssd1 vccd1 vccd1 _17189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3205 _17424_/Q vssd1 vssd1 vccd1 vccd1 hold3205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3216 _12977_/X vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _12418_/A hold812/X vssd1 vssd1 vccd1 vccd1 _16098_/D sky130_fd_sc_hd__and2_1
Xhold3227 _17376_/Q vssd1 vssd1 vccd1 vccd1 hold3227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3238 hold5883/X vssd1 vssd1 vccd1 vccd1 hold5884/A sky130_fd_sc_hd__buf_6
XFILLER_0_23_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3249 _09993_/Y vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2504 _15631_/Q vssd1 vssd1 vccd1 vccd1 hold2504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _14187_/X vssd1 vssd1 vccd1 vccd1 _17894_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07913_ hold1523/X _07918_/B _07912_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2526 _15720_/Q vssd1 vssd1 vccd1 vccd1 hold2526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08893_ _12412_/A hold892/X vssd1 vssd1 vccd1 vccd1 _16064_/D sky130_fd_sc_hd__and2_1
Xhold2537 _15817_/Q vssd1 vssd1 vccd1 vccd1 hold2537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 _15628_/Q vssd1 vssd1 vccd1 vccd1 hold2548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1803 _17885_/Q vssd1 vssd1 vccd1 vccd1 hold1803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1814 _14629_/X vssd1 vssd1 vccd1 vccd1 _18105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _17775_/Q vssd1 vssd1 vccd1 vccd1 hold2559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1825 _17908_/Q vssd1 vssd1 vccd1 vccd1 hold1825/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1836 _15178_/X vssd1 vssd1 vccd1 vccd1 _18370_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07844_ hold2248/X _07865_/B _07843_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _07844_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1847 _17910_/Q vssd1 vssd1 vccd1 vccd1 hold1847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 _14961_/X vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 _17912_/Q vssd1 vssd1 vccd1 vccd1 hold1869/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_17_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_17_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09514_ hold3860/X _10004_/B _09513_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09447_/C _09447_/D _09447_/B vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_148_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_231_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09376_ hold725/X _15483_/B _09375_/X _18458_/Q vssd1 vssd1 vccd1 vccd1 _09376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08327_ _14330_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _15211_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08189_ _14517_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5130 _16757_/Q vssd1 vssd1 vccd1 vccd1 hold5130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5141 _10525_/X vssd1 vssd1 vccd1 vccd1 _16665_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10220_ hold2953/X hold4873/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__mux2_1
Xhold5152 _16510_/Q vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5163 _09592_/X vssd1 vssd1 vccd1 vccd1 _16354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5174 _17072_/Q vssd1 vssd1 vccd1 vccd1 hold5174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5185 _11620_/X vssd1 vssd1 vccd1 vccd1 _17030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4440 _11419_/X vssd1 vssd1 vccd1 vccd1 _16963_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10151_ hold1950/X hold4639/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_6_56_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_56_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold4451 _17249_/Q vssd1 vssd1 vccd1 vccd1 hold4451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5196 _16751_/Q vssd1 vssd1 vccd1 vccd1 hold5196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4462 _13786_/X vssd1 vssd1 vccd1 vccd1 _17715_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4473 _16464_/Q vssd1 vssd1 vccd1 vccd1 hold4473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4484 _13399_/X vssd1 vssd1 vccd1 vccd1 _17586_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3750 _17433_/Q vssd1 vssd1 vccd1 vccd1 hold3750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4495 _16994_/Q vssd1 vssd1 vccd1 vccd1 hold4495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10082_ hold1183/X hold4329/X _10190_/S vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__mux2_1
Xhold3761 _12698_/X vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_332_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17210_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3772 _16998_/Q vssd1 vssd1 vccd1 vccd1 hold3772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3783 _09757_/X vssd1 vssd1 vccd1 vccd1 _16409_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3794 _10321_/X vssd1 vssd1 vccd1 vccd1 _16597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _15199_/A hold1916/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__mux2_1
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ _15121_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14890_/X sky130_fd_sc_hd__or2_1
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13841_ _17734_/Q _13847_/B _13841_/C vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16560_ _18154_/CLK _16560_/D vssd1 vssd1 vccd1 vccd1 _16560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13772_ hold2229/X hold3511/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13773_/B sky130_fd_sc_hd__mux2_1
X_10984_ hold5521/X _11210_/B _10983_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10984_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15511_ hold999/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ _12738_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _17417_/D sky130_fd_sc_hd__and2_1
X_16491_ _18364_/CLK _16491_/D vssd1 vssd1 vccd1 vccd1 _16491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _18230_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15442_ _15480_/A _15442_/B _15442_/C _15442_/D vssd1 vssd1 vccd1 vccd1 _15442_/X
+ sky130_fd_sc_hd__or4_1
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _17394_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ hold4378/X _12344_/B _11604_/X _08145_/A vssd1 vssd1 vccd1 vccd1 _11605_/X
+ sky130_fd_sc_hd__o211a_1
X_18161_ _18219_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15373_ _15490_/A1 _15365_/X _15372_/X _15490_/B1 hold5890/A vssd1 vssd1 vccd1 vccd1
+ _15373_/X sky130_fd_sc_hd__a32o_1
X_12585_ _14362_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _17371_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17112_ _17272_/CLK _17112_/D vssd1 vssd1 vccd1 vccd1 _17112_/Q sky130_fd_sc_hd__dfxtp_1
X_14324_ _15004_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11536_ hold3996/X _11726_/B _11535_/X _12975_/A vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__o211a_1
X_18092_ _18124_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14255_ hold3082/X _14272_/B _14254_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17043_ _17825_/CLK _17043_/D vssd1 vssd1 vccd1 vccd1 _17043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11467_ hold5601/X _11753_/B _11466_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13206_ _13206_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ hold3027/X hold4022/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14186_ _14758_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11398_ hold3904/X _12314_/B _11397_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11398_/X
+ sky130_fd_sc_hd__o211a_1
X_13137_ _13137_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__and2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10349_ hold2949/X hold3726/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ hold5493/X _13067_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__mux2_2
X_17945_ _18038_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ hold5010/X _12308_/B _12018_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _12019_/X
+ sky130_fd_sc_hd__o211a_1
X_17876_ _17876_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16827_ _18331_/CLK _16827_/D vssd1 vssd1 vccd1 vccd1 _16827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16758_ _18059_/CLK _16758_/D vssd1 vssd1 vccd1 vccd1 _16758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _17744_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 _15709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16689_ _18113_/CLK _16689_/D vssd1 vssd1 vccd1 vccd1 _16689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09230_ _15559_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18428_ _18428_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ hold2035/X _09164_/B _09160_/Y _15502_/A vssd1 vssd1 vccd1 vccd1 _09161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18359_ _18391_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08112_ _15517_/A hold2106/X hold240/X vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__mux2_1
X_09092_ _15099_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ _15557_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold900 hold900/A vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 hold911/A vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 hold922/A vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold933 hold933/A vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold944 hold944/A vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__clkbuf_16
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 hold966/A vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3002 _16264_/Q vssd1 vssd1 vccd1 vccd1 hold3002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 la_data_in[20] vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3013 _14107_/X vssd1 vssd1 vccd1 vccd1 _17856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _11203_/A _09994_/B vssd1 vssd1 vccd1 vccd1 _16488_/D sky130_fd_sc_hd__nor2_1
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3024 _15526_/X vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__buf_8
Xhold3035 _16236_/Q vssd1 vssd1 vccd1 vccd1 hold3035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3046 _09316_/X vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2301 _08298_/X vssd1 vssd1 vccd1 vccd1 _15782_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2312 _17877_/Q vssd1 vssd1 vccd1 vccd1 hold2312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3057 _17788_/Q vssd1 vssd1 vccd1 vccd1 hold3057/X sky130_fd_sc_hd__dlygate4sd3_1
X_08945_ hold17/X hold739/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__mux2_1
Xhold3068 _14701_/X vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2323 _18062_/Q vssd1 vssd1 vccd1 vccd1 hold2323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3079 _13048_/X vssd1 vssd1 vccd1 vccd1 _17525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 _08188_/X vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1600 _14939_/X vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2345 _17866_/Q vssd1 vssd1 vccd1 vccd1 hold2345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2356 _08034_/X vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 _14137_/X vssd1 vssd1 vccd1 vccd1 _17870_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08876_ hold113/X hold536/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__mux2_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2367 _18024_/Q vssd1 vssd1 vccd1 vccd1 hold2367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _15774_/Q vssd1 vssd1 vccd1 vccd1 hold1622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _14249_/X vssd1 vssd1 vccd1 vccd1 _17923_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 _09165_/X vssd1 vssd1 vccd1 vccd1 _16195_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1644 _18049_/Q vssd1 vssd1 vccd1 vccd1 hold1644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 _15769_/Q vssd1 vssd1 vccd1 vccd1 hold2389/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 _14207_/X vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ hold752/X hold689/X hold764/X hold732/X vssd1 vssd1 vccd1 vccd1 _14843_/A
+ sky130_fd_sc_hd__or4b_4
Xhold1666 _17968_/Q vssd1 vssd1 vccd1 vccd1 hold1666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1677 _14617_/X vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1688 _08471_/X vssd1 vssd1 vccd1 vccd1 _15864_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1699 _17792_/Q vssd1 vssd1 vccd1 vccd1 hold1699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09438_/B _16300_/Q vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09359_ hold367/A _15219_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__or3_2
XFILLER_0_34_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _13888_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _17280_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_180_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ hold1234/X hold3862/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _14774_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__nand2_1
X_11252_ hold1501/X hold4751/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10203_ _10533_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2_1
XTAP_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ _11183_/A _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__and3_1
XTAP_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4270 _13366_/X vssd1 vssd1 vccd1 vccd1 _17575_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10134_ _10542_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4281 _17266_/Q vssd1 vssd1 vccd1 vccd1 hold4281/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4292 _15323_/X vssd1 vssd1 vccd1 vccd1 _15324_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _17334_/CLK _15991_/D vssd1 vssd1 vccd1 vccd1 hold477/A sky130_fd_sc_hd__dfxtp_1
XTAP_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17730_ _17730_/CLK _17730_/D vssd1 vssd1 vccd1 vccd1 _17730_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3580 _11724_/Y vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _15211_/A _14958_/B vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or2_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ _13286_/A _10560_/A _10064_/X vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__a21oi_1
Xhold3591 _16719_/Q vssd1 vssd1 vccd1 vccd1 hold3591/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _17722_/CLK _17661_/D vssd1 vssd1 vccd1 vccd1 _17661_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2890 _15579_/Q vssd1 vssd1 vccd1 vccd1 hold2890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14873_ hold1887/X _14880_/B _14872_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14873_/X
+ sky130_fd_sc_hd__o211a_1
X_16612_ _18232_/CLK _16612_/D vssd1 vssd1 vccd1 vccd1 _16612_/Q sky130_fd_sc_hd__dfxtp_1
X_13824_ hold5681/X _13767_/A _13823_/X vssd1 vssd1 vccd1 vccd1 _13824_/Y sky130_fd_sc_hd__a21oi_1
X_17592_ _17725_/CLK _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16543_ _18131_/CLK _16543_/D vssd1 vssd1 vccd1 vccd1 _16543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ hold2262/X _16813_/Q _11159_/C vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__mux2_1
X_13755_ _13791_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_230_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ hold1121/X hold3781/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16474_ _18327_/CLK _16474_/D vssd1 vssd1 vccd1 vccd1 _16474_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ hold2299/X hold5188/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10899_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13686_ _13791_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18213_ _18213_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ _15425_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ hold3023/X _17390_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18144_ _18144_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15356_ _17339_/Q _15448_/B1 _15485_/B1 hold478/X vssd1 vssd1 vccd1 vccd1 _15356_/X
+ sky130_fd_sc_hd__a22o_1
X_12568_ hold2488/X _17367_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14307_ hold3222/X hold756/X _14306_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _14307_/X
+ sky130_fd_sc_hd__o211a_1
X_11519_ hold2985/X _16997_/Q _11711_/S vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__mux2_1
X_18075_ _18202_/CLK _18075_/D vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
X_12499_ hold2/X _12509_/A2 _12507_/A3 _12498_/X _09061_/A vssd1 vssd1 vccd1 vccd1
+ hold3/A sky130_fd_sc_hd__o311a_1
X_15287_ hold428/X _15487_/A2 _15484_/B1 hold167/X _15286_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/B sky130_fd_sc_hd__a221o_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _17904_/CLK _17026_/D vssd1 vssd1 vccd1 vccd1 _17026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14238_ _14972_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_254_wb_clk_i clkbuf_6_59_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18229_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14169_ hold1803/X _14198_/B _14168_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _14169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 _15374_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__clkbuf_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A _08934_/A vssd1 vssd1 vccd1 vccd1 _08759_/S sky130_fd_sc_hd__or2_4
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17960_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08661_ hold150/X hold699/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold700/A sky130_fd_sc_hd__mux2_1
X_17859_ _17901_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08592_ hold498/X hold907/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold908/A sky130_fd_sc_hd__mux2_1
XFILLER_0_89_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09213_ hold2401/X _09216_/B _09212_/Y _12894_/A vssd1 vssd1 vccd1 vccd1 _09213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09144_ hold944/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ hold2568/X _09119_/A2 _09074_/X _12999_/A vssd1 vssd1 vccd1 vccd1 _09075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08026_ hold2648/X _08029_/B _08025_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 hold730/A vssd1 vssd1 vccd1 vccd1 input58/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 hold752/A vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__clkbuf_4
Xhold763 input57/X vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__buf_1
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold785 hold785/A vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold796 hold796/A vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09977_ hold2691/X hold4733/X _10601_/C vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2120 _18078_/Q vssd1 vssd1 vccd1 vccd1 hold2120/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2131 _07927_/X vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2142 input69/X vssd1 vssd1 vccd1 vccd1 hold2142/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ hold292/X hold832/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__mux2_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2153 _17809_/Q vssd1 vssd1 vccd1 vccd1 hold2153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 _15619_/Q vssd1 vssd1 vccd1 vccd1 hold2164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 _18263_/Q vssd1 vssd1 vccd1 vccd1 hold1430/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2175 _08408_/X vssd1 vssd1 vccd1 vccd1 _15834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _13012_/X vssd1 vssd1 vccd1 vccd1 _17514_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2186 _16222_/Q vssd1 vssd1 vccd1 vccd1 hold2186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _18384_/Q vssd1 vssd1 vccd1 vccd1 hold1452/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2197 _17900_/Q vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ _12424_/A hold653/X vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__and2_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1463 _08312_/X vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1474 _15786_/Q vssd1 vssd1 vccd1 vccd1 hold1474/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _15640_/Q vssd1 vssd1 vccd1 vccd1 hold1485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_6_26_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _08288_/X vssd1 vssd1 vccd1 vccd1 _15777_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ hold2386/X _17114_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__mux2_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _11658_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10821_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10752_ _11136_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__or2_1
X_13540_ hold5741/X _13832_/B _13539_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13471_ hold4285/X _13886_/B _13470_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10683_ _11106_/A _10683_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12422_ _12426_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _17304_/D sky130_fd_sc_hd__and2_1
X_15210_ hold1893/X _15221_/B _15209_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _17877_/CLK _16190_/D vssd1 vssd1 vccd1 vccd1 _16190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15141_ _15195_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ _17275_/Q _12353_/B _13793_/S vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ _12234_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11304_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15072_ _15072_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12284_ hold2658/X hold4946/X _12317_/C vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14023_ hold2854/X _14040_/B _14022_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _14023_/X
+ sky130_fd_sc_hd__o211a_1
X_11235_ _12213_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ hold3591/X _11643_/A _11165_/X vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10117_ hold5407/X _10619_/B _10116_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _17293_/CLK _15974_/D vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__dfxtp_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11097_/X sky130_fd_sc_hd__or2_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17745_/CLK _17713_/D vssd1 vssd1 vccd1 vccd1 _17713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ _10603_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _16506_/D sky130_fd_sc_hd__nor2_1
X_14925_ hold2679/X _14952_/B _14924_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _14925_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17644_ _17740_/CLK _17644_/D vssd1 vssd1 vccd1 vccd1 _17644_/Q sky130_fd_sc_hd__dfxtp_1
X_14856_ _15195_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__or2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13807_ _13825_/A _13807_/B vssd1 vssd1 vccd1 vccd1 _17722_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_231_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17575_ _17607_/CLK _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14787_ hold2865/X _14774_/B _14786_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14787_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11999_ hold2156/X _17157_/Q _12302_/C vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16526_ _18224_/CLK _16526_/D vssd1 vssd1 vccd1 vccd1 _16526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13738_ hold5729/X _13817_/B _13737_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13738_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16457_ _18373_/CLK _16457_/D vssd1 vssd1 vccd1 vccd1 _16457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13669_ hold4567/X _13883_/B _13668_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15408_ hold641/X _15484_/A2 _09392_/D hold492/X vssd1 vssd1 vccd1 vccd1 _15408_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16388_ _18363_/CLK _16388_/D vssd1 vssd1 vccd1 vccd1 _16388_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_435_wb_clk_i clkbuf_6_10_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17730_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18127_ _18223_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_1
X_15339_ hold702/X _15485_/A2 _15488_/A2 hold827/X _15338_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_26_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5707 _17663_/Q vssd1 vssd1 vccd1 vccd1 hold5707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5718 _13636_/X vssd1 vssd1 vccd1 vccd1 _17665_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5729 _17731_/Q vssd1 vssd1 vccd1 vccd1 hold5729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18058_ _18058_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _09918_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17009_ _17887_/CLK _17009_/D vssd1 vssd1 vccd1 vccd1 _17009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout506 _10565_/C vssd1 vssd1 vccd1 vccd1 _10049_/C sky130_fd_sc_hd__buf_6
XFILLER_0_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout517 _10400_/S vssd1 vssd1 vccd1 vccd1 _10613_/C sky130_fd_sc_hd__clkbuf_8
X_09831_ _09843_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__or2_1
Xfanout528 _09218_/B vssd1 vssd1 vccd1 vccd1 _09216_/B sky130_fd_sc_hd__buf_4
Xfanout539 _08808_/S vssd1 vssd1 vccd1 vccd1 _08858_/S sky130_fd_sc_hd__buf_8
XFILLER_0_226_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _09954_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08713_ hold578/X hold633/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_198_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09693_ _11064_/A _09693_/B vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ _12396_/A hold839/X vssd1 vssd1 vccd1 vccd1 _15944_/D sky130_fd_sc_hd__and2_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ _12386_/A hold325/X vssd1 vssd1 vccd1 vccd1 _15911_/D sky130_fd_sc_hd__and2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_176_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18349_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09127_ hold1464/X _09177_/A2 _09126_/X _12921_/A vssd1 vssd1 vccd1 vccd1 _09127_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_105_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17301_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ hold292/X hold294/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ _15523_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__or2_1
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold571 hold97/X vssd1 vssd1 vccd1 vccd1 input6/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 hold582/A vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ hold4459/X _11762_/B _11019_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o211a_1
Xhold593 hold593/A vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _17500_/Q hold2144/X _12974_/S vssd1 vssd1 vccd1 vccd1 _12971_/X sky130_fd_sc_hd__mux2_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 _15826_/Q vssd1 vssd1 vccd1 vccd1 hold1260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14710_ _15103_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14710_/X sky130_fd_sc_hd__or2_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1271 _17779_/Q vssd1 vssd1 vccd1 vccd1 hold1271/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _14311_/X vssd1 vssd1 vccd1 vccd1 _17953_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _12213_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__or2_1
XFILLER_0_197_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1293 _15552_/X vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ _17278_/CLK _15690_/D vssd1 vssd1 vccd1 vccd1 _15690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14641_ hold2750/X _14664_/B _14640_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14641_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _13773_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__or2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ hold5188/X _11198_/B _10803_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10804_/X
+ sky130_fd_sc_hd__o211a_1
X_17360_ _17379_/CLK _17360_/D vssd1 vssd1 vccd1 vccd1 _17360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14572_ hold238/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14572_/X sky130_fd_sc_hd__and2_1
X_11784_ hold4857/X _12234_/A _11783_/X vssd1 vssd1 vccd1 vccd1 _11784_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _16311_/CLK _16311_/D vssd1 vssd1 vccd1 vccd1 _16311_/Q sky130_fd_sc_hd__dfxtp_1
X_13523_ hold2290/X hold4044/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ _18401_/CLK _17291_/D vssd1 vssd1 vccd1 vccd1 hold778/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ hold4105/X _11198_/B _10734_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _17422_/CLK _16242_/D vssd1 vssd1 vccd1 vccd1 _16242_/Q sky130_fd_sc_hd__dfxtp_1
X_10666_ hold5503/X _11156_/B _10665_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10666_/X
+ sky130_fd_sc_hd__o211a_1
X_13454_ _15842_/Q _17605_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ hold271/X hold574/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__mux2_1
X_13385_ hold2151/X hold4012/X _13826_/C vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__mux2_1
X_16173_ _17509_/CLK _16173_/D vssd1 vssd1 vccd1 vccd1 _16173_/Q sky130_fd_sc_hd__dfxtp_1
X_10597_ _18461_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _16689_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15124_ hold5980/X _15111_/B hold735/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 hold736/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput109 hold5833/X vssd1 vssd1 vccd1 vccd1 hold5834/A sky130_fd_sc_hd__buf_6
X_12336_ hold3627/X _13461_/A _12335_/X vssd1 vssd1 vccd1 vccd1 _12336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ hold246/X hold741/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold742/A sky130_fd_sc_hd__mux2_1
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12267_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _16896_/D sky130_fd_sc_hd__nor2_1
X_14006_ _14794_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__or2_1
X_12198_ _12288_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__or2_1
Xoutput80 _13193_/A vssd1 vssd1 vccd1 vccd1 output80/X sky130_fd_sc_hd__buf_6
Xoutput91 _13273_/A vssd1 vssd1 vccd1 vccd1 output91/X sky130_fd_sc_hd__buf_6
XFILLER_0_208_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11149_ _11158_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _16873_/D sky130_fd_sc_hd__nor2_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ _17304_/CLK _15957_/D vssd1 vssd1 vccd1 vccd1 hold785/A sky130_fd_sc_hd__dfxtp_1
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ hold525/X _14910_/B vssd1 vssd1 vccd1 vccd1 hold526/A sky130_fd_sc_hd__or2_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15888_ _17334_/CLK _15888_/D vssd1 vssd1 vccd1 vccd1 hold725/A sky130_fd_sc_hd__dfxtp_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17627_ _17721_/CLK _17627_/D vssd1 vssd1 vccd1 vccd1 _17627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ hold1718/X _14826_/B _14838_/X _14839_/C1 vssd1 vssd1 vccd1 vccd1 _14839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_231_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08360_ _15529_/A hold2596/X hold134/X vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17558_ _17718_/CLK _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _18362_/CLK _16509_/D vssd1 vssd1 vccd1 vccd1 _16509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08291_ _14116_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08291_/X sky130_fd_sc_hd__or2_1
X_17489_ _17491_/CLK _17489_/D vssd1 vssd1 vccd1 vccd1 _17489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5504 _10666_/X vssd1 vssd1 vccd1 vccd1 _16712_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5515 _16882_/Q vssd1 vssd1 vccd1 vccd1 hold5515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5526 _11485_/X vssd1 vssd1 vccd1 vccd1 _16985_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5537 _16947_/Q vssd1 vssd1 vccd1 vccd1 hold5537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4803 _16603_/Q vssd1 vssd1 vccd1 vccd1 hold4803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5548 _11584_/X vssd1 vssd1 vccd1 vccd1 _17018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4814 _10510_/X vssd1 vssd1 vccd1 vccd1 _16660_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5559 _16814_/Q vssd1 vssd1 vccd1 vccd1 hold5559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4825 _16756_/Q vssd1 vssd1 vccd1 vccd1 hold4825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4836 _10183_/X vssd1 vssd1 vccd1 vccd1 _16551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4847 _16650_/Q vssd1 vssd1 vccd1 vccd1 hold4847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4858 _11784_/Y vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout303 _09918_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__buf_4
Xhold4869 _16690_/Q vssd1 vssd1 vccd1 vccd1 hold4869/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout314 _11094_/A vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__buf_4
Xfanout325 _09564_/A vssd1 vssd1 vccd1 vccd1 _10488_/A sky130_fd_sc_hd__buf_4
XFILLER_0_226_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout336 _12500_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__buf_4
Xfanout347 _08932_/S vssd1 vssd1 vccd1 vccd1 _08928_/S sky130_fd_sc_hd__buf_6
X_09814_ hold3898/X _10004_/B _09813_/X _15234_/C1 vssd1 vssd1 vccd1 vccd1 _09814_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout358 _15560_/A2 vssd1 vssd1 vccd1 vccd1 _15547_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout369 hold394/X vssd1 vssd1 vccd1 vccd1 _15071_/S sky130_fd_sc_hd__buf_8
XFILLER_0_241_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ hold3858/X _10007_/B _09744_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09745_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ hold5679/X _10070_/B _09675_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08627_ hold118/X hold458/X _08627_/S vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08558_ hold454/X hold840/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold841/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_357_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08489_ hold2288/X _08486_/B _08488_/Y _08381_/A vssd1 vssd1 vccd1 vccd1 _08489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ hold1147/X _16664_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ hold1937/X hold3956/X _10997_/S vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _17572_/Q _17106_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__mux2_1
X_10382_ hold2176/X _16618_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ hold5405/X _13862_/B _12120_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ hold5599/X _12052_/A2 _12051_/X _08127_/A vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o211a_1
Xhold390 input61/X vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11003_ hold2733/X hold4240/X _11192_/C vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_73_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17372_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _18061_/CLK _16860_/D vssd1 vssd1 vccd1 vccd1 _16860_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout870 fanout873/X vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__clkbuf_8
X_15811_ _17658_/CLK _15811_/D vssd1 vssd1 vccd1 vccd1 _15811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 hold1107/X vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__clkbuf_16
X_16791_ _18230_/CLK _16791_/D vssd1 vssd1 vccd1 vccd1 _16791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout892 hold926/X vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__buf_12
XFILLER_0_204_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15742_ _17745_/CLK _15742_/D vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12990_/A _12954_/B vssd1 vssd1 vccd1 vccd1 _17494_/D sky130_fd_sc_hd__and2_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 _16263_/Q vssd1 vssd1 vccd1 vccd1 hold1090/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18461_/A vssd1 vssd1 vccd1 vccd1 _18461_/X sky130_fd_sc_hd__buf_1
X_11905_ hold5160/X _13798_/A2 _11904_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15673_ _17199_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12990_/A _12885_/B vssd1 vssd1 vccd1 vccd1 _17471_/D sky130_fd_sc_hd__and2_1
XFILLER_0_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _17413_/CLK _17412_/D vssd1 vssd1 vccd1 vccd1 _17412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _15233_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__or2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18394_/CLK hold974/X vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
X_11836_ hold5391/X _12031_/A2 _11835_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17343_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _17343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14555_ _18459_/Q _14555_/B _14555_/C vssd1 vssd1 vccd1 vccd1 _14573_/B sky130_fd_sc_hd__and3_4
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _12367_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _17079_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13506_ _13698_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__or2_1
X_10718_ hold2842/X hold4676/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__mux2_1
X_17274_ _17274_/CLK _17274_/D vssd1 vssd1 vccd1 vccd1 _17274_/Q sky130_fd_sc_hd__dfxtp_1
X_14486_ hold2937/X _14487_/B _14485_/Y _14366_/A vssd1 vssd1 vccd1 vccd1 _14486_/X
+ sky130_fd_sc_hd__o211a_1
X_11698_ hold4368/X _11801_/B _11697_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11698_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16225_ _18432_/CLK _16225_/D vssd1 vssd1 vccd1 vccd1 _16225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _13734_/A _13437_/B vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10649_ _16707_/Q _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__and3_1
XFILLER_0_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16156_ _17509_/CLK _16156_/D vssd1 vssd1 vccd1 vccd1 _16156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13368_ _13776_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15541_/A _15111_/B vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ _13864_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _17263_/D sky130_fd_sc_hd__nor2_1
X_16087_ _16087_/CLK _16087_/D vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__dfxtp_1
X_13299_ _13298_/X _16930_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__mux2_1
Xhold3409 _09601_/X vssd1 vssd1 vccd1 vccd1 _16357_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15038_ _15454_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2708 _14155_/X vssd1 vssd1 vccd1 vccd1 _17879_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2719 _15651_/Q vssd1 vssd1 vccd1 vccd1 hold2719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ hold2872/X _07865_/B _07859_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _07860_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07791_ hold391/X vssd1 vssd1 vccd1 vccd1 _14555_/C sky130_fd_sc_hd__inv_2
XFILLER_0_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16989_ _17890_/CLK _16989_/D vssd1 vssd1 vccd1 vccd1 _16989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ hold3147/X _13142_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09531_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09461_ _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__and3_1
XFILLER_0_8_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ hold3019/X _08440_/A2 _08411_/X _13672_/C1 vssd1 vssd1 vccd1 vccd1 _08412_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09392_/A _09392_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09392_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_450_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17160_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08343_ _08349_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__and2_1
XFILLER_0_175_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08274_ _15553_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6002 _18357_/Q vssd1 vssd1 vccd1 vccd1 hold6002/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6013 data_in[5] vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6024 _09443_/Y vssd1 vssd1 vccd1 vccd1 _16307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6035 _18400_/Q vssd1 vssd1 vccd1 vccd1 hold6035/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6046 _16521_/Q vssd1 vssd1 vccd1 vccd1 hold6046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5301 _10678_/X vssd1 vssd1 vccd1 vccd1 _16716_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5312 _16621_/Q vssd1 vssd1 vccd1 vccd1 hold5312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5323 _09940_/X vssd1 vssd1 vccd1 vccd1 _16470_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5334 _17037_/Q vssd1 vssd1 vccd1 vccd1 hold5334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5345 _10105_/X vssd1 vssd1 vccd1 vccd1 _16525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4600 _10581_/Y vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4611 _10068_/Y vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5356 _17230_/Q vssd1 vssd1 vccd1 vccd1 hold5356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4622 _10626_/Y vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5367 _11938_/X vssd1 vssd1 vccd1 vccd1 _17136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4633 _11187_/Y vssd1 vssd1 vccd1 vccd1 _11188_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_46_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_46_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold5378 _11353_/X vssd1 vssd1 vccd1 vccd1 _16941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4644 _13818_/Y vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5389 _17231_/Q vssd1 vssd1 vccd1 vccd1 hold5389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4655 hold6045/X vssd1 vssd1 vccd1 vccd1 hold4655/X sky130_fd_sc_hd__buf_1
Xhold3910 _16969_/Q vssd1 vssd1 vccd1 vccd1 hold3910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3921 _10252_/X vssd1 vssd1 vccd1 vccd1 _16574_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4666 _16717_/Q vssd1 vssd1 vccd1 vccd1 hold4666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4677 _11199_/Y vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3932 _16968_/Q vssd1 vssd1 vccd1 vccd1 hold3932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3943 _13327_/X vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4688 _10587_/Y vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3954 _16636_/Q vssd1 vssd1 vccd1 vccd1 hold3954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4699 _16718_/Q vssd1 vssd1 vccd1 vccd1 hold4699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3965 _09988_/X vssd1 vssd1 vccd1 vccd1 _16486_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3976 _16463_/Q vssd1 vssd1 vccd1 vccd1 hold3976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3987 _09820_/X vssd1 vssd1 vccd1 vccd1 _16430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout155 _12986_/S vssd1 vssd1 vccd1 vccd1 _12998_/S sky130_fd_sc_hd__buf_6
XFILLER_0_227_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout166 _13817_/B vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__buf_4
Xhold3998 _17033_/Q vssd1 vssd1 vccd1 vccd1 hold3998/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout177 _11747_/B vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__clkbuf_8
Xfanout188 _12347_/B vssd1 vssd1 vccd1 vccd1 _13868_/B sky130_fd_sc_hd__buf_4
Xfanout199 _11210_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__buf_4
X_07989_ hold1369/X _07991_/A2 _07988_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _07989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09728_ hold741/X hold4481/X _09824_/S vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_236_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09659_ _18288_/Q hold3631/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ hold2361/X _17401_/Q _12772_/S vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ hold2312/X _17031_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ hold331/X _14502_/B vssd1 vssd1 vccd1 vccd1 hold332/A sky130_fd_sc_hd__or2_1
XFILLER_0_167_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ hold2763/X hold5246/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _11100_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11483_ hold1561/X hold5457/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__mux2_1
X_14271_ hold1904/X _14272_/B _14270_/Y _13917_/A vssd1 vssd1 vccd1 vccd1 _14271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16010_ _18399_/CLK _16010_/D vssd1 vssd1 vccd1 vccd1 hold609/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10434_ _10533_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__or2_1
X_13222_ _13222_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13153_ _13153_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__and2_1
X_10365_ _11097_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ hold2548/X hold4915/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084_ hold3732/X _13083_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_2
X_17961_ _18200_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5890 hold5890/A vssd1 vssd1 vccd1 vccd1 hold5890/X sky130_fd_sc_hd__clkbuf_4
X_10296_ _10524_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10296_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12035_ hold2656/X _17169_/Q _12251_/S vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__mux2_1
X_16912_ _17886_/CLK _16912_/D vssd1 vssd1 vccd1 vccd1 _16912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17892_ _17892_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_1
X_16843_ _18044_/CLK _16843_/D vssd1 vssd1 vccd1 vccd1 _16843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16774_ _17975_/CLK _16774_/D vssd1 vssd1 vccd1 vccd1 _16774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_279_wb_clk_i clkbuf_6_50_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13986_ _14774_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _17728_/CLK _15725_/D vssd1 vssd1 vccd1 vccd1 _15725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ hold2049/X _17490_/Q _12997_/S vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_208_wb_clk_i clkbuf_6_55_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18444_ _18445_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15656_ _17164_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ hold1423/X hold3224/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14607_ hold2971/X _14610_/B _14606_/Y _14827_/C1 vssd1 vssd1 vccd1 vccd1 _14607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18375_ _18375_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ hold1115/X hold4672/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15587_ _17899_/CLK _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
X_12799_ hold2527/X hold3217/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ _17326_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 _17326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14538_ hold2244/X _14541_/B _14537_/Y _14538_/C1 vssd1 vssd1 vccd1 vccd1 _14538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17257_ _17257_/CLK _17257_/D vssd1 vssd1 vccd1 vccd1 _17257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14469_ _14988_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14469_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16208_ _18435_/CLK _16208_/D vssd1 vssd1 vccd1 vccd1 _16208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ _17188_/CLK _17188_/D vssd1 vssd1 vccd1 vccd1 _17188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16139_ _17314_/CLK _16139_/D vssd1 vssd1 vccd1 vccd1 hold637/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3206 _12743_/X vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3217 _17444_/Q vssd1 vssd1 vccd1 vccd1 hold3217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08961_ hold454/X hold811/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold812/A sky130_fd_sc_hd__mux2_1
Xhold3228 _12599_/X vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3239 _09394_/X vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2505 _07977_/X vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 _18177_/Q vssd1 vssd1 vccd1 vccd1 hold2516/X sky130_fd_sc_hd__dlygate4sd3_1
X_07912_ _14529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07912_/X sky130_fd_sc_hd__or2_1
Xhold2527 _16212_/Q vssd1 vssd1 vccd1 vccd1 hold2527/X sky130_fd_sc_hd__dlygate4sd3_1
X_08892_ hold361/X hold891/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold892/A sky130_fd_sc_hd__mux2_1
Xhold2538 _15636_/Q vssd1 vssd1 vccd1 vccd1 hold2538/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 _14169_/X vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 _07971_/X vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 _16298_/Q vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07843_ _15521_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07843_/X sky130_fd_sc_hd__or2_1
Xhold1826 _14215_/X vssd1 vssd1 vccd1 vccd1 _17908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1837 _17994_/Q vssd1 vssd1 vccd1 vccd1 hold1837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1848 _14221_/X vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _18178_/Q vssd1 vssd1 vccd1 vccd1 hold1859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _09987_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__and3_1
XFILLER_0_56_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _15480_/A _09375_/B _09375_/C _09375_/D vssd1 vssd1 vccd1 vccd1 _09375_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08326_ hold2047/X _08336_/A2 _08325_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ hold1605/X _08263_/A2 _08256_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _08257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08188_ hold2333/X _08209_/B _08187_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5120 _16956_/Q vssd1 vssd1 vccd1 vccd1 hold5120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5131 _10705_/X vssd1 vssd1 vccd1 vccd1 _16725_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5142 _16791_/Q vssd1 vssd1 vccd1 vccd1 hold5142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5153 _09964_/X vssd1 vssd1 vccd1 vccd1 _16478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5164 _16890_/Q vssd1 vssd1 vccd1 vccd1 hold5164/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5175 _11650_/X vssd1 vssd1 vccd1 vccd1 _17040_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4430 _11116_/X vssd1 vssd1 vccd1 vccd1 _16862_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10150_ hold3902/X _10628_/B _10149_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10150_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4441 _17651_/Q vssd1 vssd1 vccd1 vccd1 hold4441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5186 _17163_/Q vssd1 vssd1 vccd1 vccd1 hold5186/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4452 _12181_/X vssd1 vssd1 vccd1 vccd1 _17217_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5197 _10687_/X vssd1 vssd1 vccd1 vccd1 _16719_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4463 _17091_/Q vssd1 vssd1 vccd1 vccd1 hold4463/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4474 _09826_/X vssd1 vssd1 vccd1 vccd1 _16432_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3740 _17586_/Q vssd1 vssd1 vccd1 vccd1 hold3740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4485 _17175_/Q vssd1 vssd1 vccd1 vccd1 hold4485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ hold4775/X _10565_/B _10080_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _10081_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3751 _12770_/X vssd1 vssd1 vccd1 vccd1 _12771_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4496 _11416_/X vssd1 vssd1 vccd1 vccd1 _16962_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3762 _16966_/Q vssd1 vssd1 vccd1 vccd1 hold3762/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3773 _11428_/X vssd1 vssd1 vccd1 vccd1 _16966_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3784 _17061_/Q vssd1 vssd1 vccd1 vccd1 hold3784/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3795 _17400_/Q vssd1 vssd1 vccd1 vccd1 hold3795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13840_ _13873_/A _13840_/B vssd1 vssd1 vccd1 vccd1 _17733_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_372_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ hold4565/X _13856_/B _13770_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10983_ _11658_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_301_wb_clk_i clkbuf_6_38_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17860_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ hold1432/X _15507_/Y _15509_/X _12870_/A vssd1 vssd1 vccd1 vccd1 _15510_/X
+ sky130_fd_sc_hd__o211a_1
X_12722_ hold3372/X _12721_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__mux2_1
X_16490_ _18273_/CLK _16490_/D vssd1 vssd1 vccd1 vccd1 _16490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15441_ hold788/X _15451_/A2 _09386_/D hold801/X _15436_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/D sky130_fd_sc_hd__a221o_1
X_12653_ hold3701/X _12652_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__mux2_1
X_18160_ _18222_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
X_11604_ _12057_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__or2_1
X_15372_ _15489_/A _15372_/B _15372_/C _15372_/D vssd1 vssd1 vccd1 vccd1 _15372_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_182_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12584_ hold3175/X _12583_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17111_ _17207_/CLK _17111_/D vssd1 vssd1 vccd1 vccd1 _17111_/Q sky130_fd_sc_hd__dfxtp_1
X_14323_ hold2190/X _14326_/B _14322_/Y _14388_/A vssd1 vssd1 vccd1 vccd1 _14323_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18091_ _18123_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11535_ _11631_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _17888_/CLK _17042_/D vssd1 vssd1 vccd1 vccd1 _17042_/Q sky130_fd_sc_hd__dfxtp_1
X_14254_ _14988_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ _11658_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _13204_/X hold3581/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__mux2_1
X_10417_ hold4954/X _10631_/B _10416_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11397_ _12219_/A _11397_/B vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14185_ hold1626/X _14202_/B _14184_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _13129_/X _13135_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17535_/D sky130_fd_sc_hd__o21a_1
X_10348_ hold5136/X _11095_/A2 _10347_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ hold5170/X _10571_/B _10278_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10279_/X
+ sky130_fd_sc_hd__o211a_1
X_17944_ _18012_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13066_/X _16901_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ _12213_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_206_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17875_ _17875_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16826_ _18032_/CLK _16826_/D vssd1 vssd1 vccd1 vccd1 _16826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16757_ _18054_/CLK _16757_/D vssd1 vssd1 vccd1 vccd1 _16757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13969_ hold2961/X _13995_/A2 _13968_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _13969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15708_ _17276_/CLK hold242/X vssd1 vssd1 vccd1 vccd1 _15708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ _18208_/CLK _16688_/D vssd1 vssd1 vccd1 vccd1 _16688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _17272_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_1
X_18427_ _18427_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _15543_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09160_/Y sky130_fd_sc_hd__nand2_1
X_18358_ _18390_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__and2_1
X_17309_ _17523_/CLK _17309_/D vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09091_ hold2455/X _09106_/B _09090_/X _12960_/A vssd1 vssd1 vccd1 vccd1 _09091_/X
+ sky130_fd_sc_hd__o211a_1
X_18289_ _18353_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ hold2282/X _08033_/B _08041_/X _08385_/A vssd1 vssd1 vccd1 vccd1 _08042_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold901 hold901/A vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 hold912/A vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/A vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold934 hold934/A vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold945 hold945/A vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 hold967/A vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3003 _09308_/X vssd1 vssd1 vccd1 vccd1 _16264_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 input49/A sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _13094_/A _09918_/A _09992_/X vssd1 vssd1 vccd1 vccd1 _09993_/Y sky130_fd_sc_hd__a21oi_1
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3014 _17756_/Q vssd1 vssd1 vccd1 vccd1 hold3014/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3025 _18193_/Q vssd1 vssd1 vccd1 vccd1 hold3025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3036 _18034_/Q vssd1 vssd1 vccd1 vccd1 hold3036/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3047 _18104_/Q vssd1 vssd1 vccd1 vccd1 hold3047/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2302 _15606_/Q vssd1 vssd1 vccd1 vccd1 hold2302/X sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ _15264_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _16089_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2313 _14151_/X vssd1 vssd1 vccd1 vccd1 _17877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3058 _13967_/X vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 _18008_/Q vssd1 vssd1 vccd1 vccd1 hold3069/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 _14536_/X vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2335 _15624_/Q vssd1 vssd1 vccd1 vccd1 hold2335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 _18294_/Q vssd1 vssd1 vccd1 vccd1 hold1601/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2346 _14129_/X vssd1 vssd1 vccd1 vccd1 _17866_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1612 _18214_/Q vssd1 vssd1 vccd1 vccd1 hold1612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 _15674_/Q vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__dlygate4sd3_1
X_08875_ _12386_/A hold474/X vssd1 vssd1 vccd1 vccd1 _16055_/D sky130_fd_sc_hd__and2_1
Xhold1623 _08279_/X vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2368 _14458_/X vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1634 _18059_/Q vssd1 vssd1 vccd1 vccd1 hold1634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 _15816_/Q vssd1 vssd1 vccd1 vccd1 hold2379/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1645 _14510_/X vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ _07826_/A _13048_/A vssd1 vssd1 vccd1 vccd1 _07826_/X sky130_fd_sc_hd__and2_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1656 _17818_/Q vssd1 vssd1 vccd1 vccd1 hold1656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1667 _14341_/X vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1678 _18269_/Q vssd1 vssd1 vccd1 vccd1 hold1678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1689 _18331_/Q vssd1 vssd1 vccd1 vccd1 hold1689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09427_ _07804_/A _09472_/B _15344_/A _09426_/X vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09358_ _09366_/A _09363_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09358_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08309_ _15533_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08309_/X sky130_fd_sc_hd__or2_1
X_09289_ hold999/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11320_ hold3525/X _11584_/A2 _11319_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ hold4069/X _11729_/B _11250_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ hold3090/X hold5064/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11182_ _11194_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _16884_/D sky130_fd_sc_hd__nor2_1
XTAP_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4260 _13684_/X vssd1 vssd1 vccd1 vccd1 _17681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_235_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ hold2884/X hold3549/X _10613_/C vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__mux2_1
Xhold4271 hold5840/X vssd1 vssd1 vccd1 vccd1 hold4271/X sky130_fd_sc_hd__buf_4
XTAP_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15990_ _17335_/CLK _15990_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4282 _12232_/X vssd1 vssd1 vccd1 vccd1 _17234_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4293 _17024_/Q vssd1 vssd1 vccd1 vccd1 hold4293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3570 _12303_/Y vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10064_ _16512_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__and3_1
Xhold3581 _16534_/Q vssd1 vssd1 vccd1 vccd1 hold3581/X sky130_fd_sc_hd__buf_1
X_14941_ hold1581/X _14952_/B _14940_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14941_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3592 _11166_/Y vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _18447_/CLK _17660_/D vssd1 vssd1 vccd1 vccd1 _17660_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2880 _15563_/Q vssd1 vssd1 vccd1 vccd1 hold2880/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _15211_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__or2_1
Xhold2891 _07868_/X vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16611_ _18231_/CLK _16611_/D vssd1 vssd1 vccd1 vccd1 _16611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13823_ _17728_/Q _13832_/B _13826_/C vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__and3_1
X_17591_ _17623_/CLK _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16542_ _18182_/CLK _16542_/D vssd1 vssd1 vccd1 vccd1 _16542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13754_ hold2945/X _17705_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10966_ hold3535/X _11156_/B _10965_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _10966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12705_ _12768_/A _12705_/B vssd1 vssd1 vccd1 vccd1 _17411_/D sky130_fd_sc_hd__and2_1
X_16473_ _18384_/CLK _16473_/D vssd1 vssd1 vccd1 vccd1 _16473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13685_ hold1605/X hold3458/X _13874_/C vssd1 vssd1 vccd1 vccd1 _13686_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10897_ hold3841/X _11095_/A2 _10896_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18212_ _18212_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _15454_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__and2_1
XFILLER_0_122_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12636_ _12810_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _17388_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ _18143_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ hold668/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12567_ _12960_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _17365_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _15201_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18074_ _18265_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11518_ hold5342/X _12317_/B _11517_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11518_/X
+ sky130_fd_sc_hd__o211a_1
X_15286_ _17332_/Q _15448_/B1 _15485_/B1 hold592/X vssd1 vssd1 vccd1 vccd1 _15286_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12498_ _17342_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__or2_1
Xhold208 hold1/X vssd1 vssd1 vccd1 vccd1 input23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17025_ _17871_/CLK _17025_/D vssd1 vssd1 vccd1 vccd1 _17025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14237_ hold1442/X _14266_/B _14236_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14237_/X
+ sky130_fd_sc_hd__o211a_1
X_11449_ hold5292/X _11732_/B _11448_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ _14972_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_221_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13199_/A1 _13117_/X _13118_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_294_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ hold1391/X _14094_/B _14098_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _18226_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_223_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18215_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08660_ _12412_/A hold910/X vssd1 vssd1 vccd1 vccd1 _15952_/D sky130_fd_sc_hd__and2_1
X_17858_ _17858_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16809_ _18010_/CLK _16809_/D vssd1 vssd1 vccd1 vccd1 _16809_/Q sky130_fd_sc_hd__dfxtp_1
X_08591_ _15304_/A hold829/X vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17789_ _17885_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_232_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09212_ _15541_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ hold3039/X _09164_/B _09142_/X _12912_/A vssd1 vssd1 vccd1 vccd1 _09143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ _15515_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08025_ _15539_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 hold720/A vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 input58/X vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 hold764/A vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__buf_2
XFILLER_0_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold775 hold775/A vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold797/A vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ hold5699/X _10468_/A2 _09975_/X _09976_/C1 vssd1 vssd1 vccd1 vccd1 _09976_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2110 _14568_/X vssd1 vssd1 vccd1 vccd1 hold2110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2121 _14570_/X vssd1 vssd1 vccd1 vccd1 hold2121/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2132 _17887_/Q vssd1 vssd1 vccd1 vccd1 hold2132/X sky130_fd_sc_hd__dlygate4sd3_1
X_08927_ _15414_/A hold357/X vssd1 vssd1 vccd1 vccd1 _16081_/D sky130_fd_sc_hd__and2_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2143 _12513_/X vssd1 vssd1 vccd1 vccd1 _12970_/S sky130_fd_sc_hd__buf_4
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2154 _14011_/X vssd1 vssd1 vccd1 vccd1 _17809_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _07953_/X vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 _17806_/Q vssd1 vssd1 vccd1 vccd1 hold1420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 _14957_/X vssd1 vssd1 vccd1 vccd1 _18263_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2176 _18174_/Q vssd1 vssd1 vccd1 vccd1 hold2176/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1442 _17917_/Q vssd1 vssd1 vccd1 vccd1 hold1442/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ hold145/X hold652/X _08858_/S vssd1 vssd1 vccd1 vccd1 hold653/A sky130_fd_sc_hd__mux2_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2187 _09221_/X vssd1 vssd1 vccd1 vccd1 _16222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _15208_/X vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2198 _14199_/X vssd1 vssd1 vccd1 vccd1 _17900_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 _16176_/Q vssd1 vssd1 vccd1 vccd1 hold1464/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1475 _08306_/X vssd1 vssd1 vccd1 vccd1 _15786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07809_ _18457_/Q _18458_/Q vssd1 vssd1 vccd1 vccd1 _07809_/X sky130_fd_sc_hd__or2_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1486 _07998_/X vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1497 _18279_/Q vssd1 vssd1 vccd1 vccd1 hold1497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08789_ hold292/X _16015_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__mux2_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ hold2449/X hold4453/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_98_wb_clk_i clkbuf_6_22_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ hold1958/X _16741_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _13779_/A _13470_/B vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_6_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17508_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10682_ hold3185/X hold4699/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10683_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ hold353/X hold788/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_6_5_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_15140_ hold3029/X _15167_/B _15139_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15140_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12352_ _13873_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _17274_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _17771_/Q hold4857/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__mux2_1
X_15071_ _15233_/A hold2973/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__mux2_1
X_12283_ hold4411/X _13877_/B _12282_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12283_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _15529_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11234_ hold1544/X hold5106/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _16879_/Q _11738_/B _11168_/C vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__and3_1
XTAP_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4090 _13702_/X vssd1 vssd1 vccd1 vccd1 _17687_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _10524_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__or2_1
XTAP_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15973_ _17327_/CLK _15973_/D vssd1 vssd1 vccd1 vccd1 _15973_/Q sky130_fd_sc_hd__dfxtp_1
X_11096_ hold2542/X _16856_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__mux2_1
XTAP_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ _13238_/A _09954_/A _10046_/X vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__a21oi_1
X_14924_ _15193_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__or2_1
X_17712_ _17712_/CLK _17712_/D vssd1 vssd1 vccd1 vccd1 _17712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__buf_1
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ hold1612/X _14882_/B _14854_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14855_/X
+ sky130_fd_sc_hd__o211a_1
X_17643_ _17707_/CLK _17643_/D vssd1 vssd1 vccd1 vccd1 _17643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13806_ hold3565/X _13623_/A _13805_/X vssd1 vssd1 vccd1 vccd1 _13806_/Y sky130_fd_sc_hd__a21oi_1
X_17574_ _17734_/CLK _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14786_ _15233_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14786_/X sky130_fd_sc_hd__or2_1
X_11998_ hold4253/X _12353_/B _11997_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__o211a_1
X_16525_ _18113_/CLK _16525_/D vssd1 vssd1 vccd1 vccd1 _16525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13737_ _13767_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__or2_1
X_10949_ hold3069/X hold4283/X _11147_/C vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16456_ _18367_/CLK _16456_/D vssd1 vssd1 vccd1 vccd1 _16456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13668_ _13788_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15407_ _17316_/Q _15487_/A2 _15484_/B1 hold234/X _15406_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12619_ hold2054/X hold3310/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__mux2_1
X_16387_ _18266_/CLK _16387_/D vssd1 vssd1 vccd1 vccd1 _16387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13599_ _13779_/A _13599_/B vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _18152_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ hold643/X _15484_/A2 _09392_/D hold670/X vssd1 vssd1 vccd1 vccd1 _15338_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5708 _13534_/X vssd1 vssd1 vccd1 vccd1 _17631_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5719 _17677_/Q vssd1 vssd1 vccd1 vccd1 hold5719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18057_ _18226_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15269_ hold430/X _15485_/A2 _09392_/C hold768/X _15268_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_223_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _17886_/CLK _17008_/D vssd1 vssd1 vccd1 vccd1 _17008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_404_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17852_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout507 _10565_/C vssd1 vssd1 vccd1 vccd1 _10571_/C sky130_fd_sc_hd__clkbuf_8
X_09830_ hold3033/X hold4535/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout518 _10025_/C vssd1 vssd1 vccd1 vccd1 _10400_/S sky130_fd_sc_hd__buf_8
XFILLER_0_1_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout529 _09178_/Y vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__buf_4
X_09761_ _18322_/Q hold3635/X _10565_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08712_ _15324_/A hold461/X vssd1 vssd1 vccd1 vccd1 _15977_/D sky130_fd_sc_hd__and2_1
XFILLER_0_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09692_ hold2544/X _16388_/Q _09824_/S vssd1 vssd1 vccd1 vccd1 _09693_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08643_ hold607/X hold838/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold839/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08574_ hold228/X hold324/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09126_ _15509_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _12438_/A hold141/X vssd1 vssd1 vccd1 vccd1 _16145_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ hold2156/X _08029_/B _08007_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _08008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_145_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_198_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold550 hold550/A vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 input6/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold583 hold583/A vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 hold70/X vssd1 vssd1 vccd1 vccd1 input34/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ hold1212/X hold4749/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__mux2_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _16164_/Q _17501_/Q _12970_/S vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_231_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 _08254_/X vssd1 vssd1 vccd1 vccd1 hold1250/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 _18432_/Q vssd1 vssd1 vccd1 vccd1 hold1261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ hold2227/X hold5072/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_197_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _13949_/X vssd1 vssd1 vccd1 vccd1 _17779_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1283 _18275_/Q vssd1 vssd1 vccd1 vccd1 hold1283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _15626_/Q vssd1 vssd1 vccd1 vccd1 hold1294/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14910_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ hold2168/X hold3611/X _13868_/C vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__mux2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10803_ _11103_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14571_ _14910_/A _14557_/Y hold2121/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14571_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11783_ _17085_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _11783_/X sky130_fd_sc_hd__and3_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16310_ _16311_/CLK _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/Q sky130_fd_sc_hd__dfxtp_1
X_13522_ hold4129/X _13802_/B _13521_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _13522_/X
+ sky130_fd_sc_hd__o211a_1
X_17290_ _18415_/CLK _17290_/D vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__dfxtp_1
X_10734_ _11103_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16241_ _17422_/CLK _16241_/D vssd1 vssd1 vccd1 vccd1 _16241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13453_ hold4545/X _13856_/B _13452_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10665_ _11136_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12404_ _12404_/A hold869/X vssd1 vssd1 vccd1 vccd1 _17295_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ _17509_/CLK _16172_/D vssd1 vssd1 vccd1 vccd1 _16172_/Q sky130_fd_sc_hd__dfxtp_1
X_13384_ hold5499/X _12353_/B _13383_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _13384_/X
+ sky130_fd_sc_hd__o211a_1
X_10596_ hold4725/X _10524_/A _10595_/X vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ hold719/X hold734/X vssd1 vssd1 vccd1 vccd1 hold735/A sky130_fd_sc_hd__or2_1
XFILLER_0_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12335_ _12335_/A _12374_/B _13556_/S vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ _15058_/A hold472/X vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12266_ hold2166/X _17246_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ hold1420/X _14038_/B _14004_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _14005_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11217_ hold4707/X _11121_/A _11216_/X vssd1 vssd1 vccd1 vccd1 _11217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12197_ hold2130/X hold4913/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__mux2_1
Xoutput81 _13201_/A vssd1 vssd1 vccd1 vccd1 output81/X sky130_fd_sc_hd__buf_6
Xoutput92 _13281_/A vssd1 vssd1 vccd1 vccd1 output92/X sky130_fd_sc_hd__buf_6
XFILLER_0_235_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11148_ hold3758/X _11052_/A _11147_/X vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15956_ _17303_/CLK _15956_/D vssd1 vssd1 vccd1 vccd1 hold769/A sky130_fd_sc_hd__dfxtp_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _11082_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__or2_1
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ hold940/X _14896_/Y _14906_/X _15394_/A vssd1 vssd1 vccd1 vccd1 hold941/A
+ sky130_fd_sc_hd__o211a_1
X_15887_ _18423_/CLK _15887_/D vssd1 vssd1 vccd1 vccd1 hold790/A sky130_fd_sc_hd__dfxtp_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17626_ _17658_/CLK _17626_/D vssd1 vssd1 vccd1 vccd1 _17626_/Q sky130_fd_sc_hd__dfxtp_1
X_14838_ _15231_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ _18131_/CLK _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
X_14769_ hold2852/X _14772_/B _14768_/Y _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14769_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16508_ _18387_/CLK _16508_/D vssd1 vssd1 vccd1 vccd1 _16508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08290_ hold2723/X _08323_/B _08289_/X _08369_/A vssd1 vssd1 vccd1 vccd1 _08290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17488_ _17491_/CLK _17488_/D vssd1 vssd1 vccd1 vccd1 _17488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16439_ _18382_/CLK _16439_/D vssd1 vssd1 vccd1 vccd1 _16439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5505 _16986_/Q vssd1 vssd1 vccd1 vccd1 hold5505/X sky130_fd_sc_hd__dlygate4sd3_1
X_18109_ _18178_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5516 _11080_/X vssd1 vssd1 vccd1 vccd1 _16850_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5527 _16498_/Q vssd1 vssd1 vccd1 vccd1 hold5527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5538 _11275_/X vssd1 vssd1 vccd1 vccd1 _16915_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4804 _10243_/X vssd1 vssd1 vccd1 vccd1 _16571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_6_36_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_36_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
Xhold5549 _16766_/Q vssd1 vssd1 vccd1 vccd1 hold5549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4815 _16918_/Q vssd1 vssd1 vccd1 vccd1 hold4815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4826 _10702_/X vssd1 vssd1 vccd1 vccd1 _16724_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4837 _16436_/Q vssd1 vssd1 vccd1 vccd1 hold4837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4848 _10384_/X vssd1 vssd1 vccd1 vccd1 _16618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4859 _16618_/Q vssd1 vssd1 vccd1 vccd1 hold4859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout304 _11061_/A vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__buf_4
Xfanout315 _11094_/A vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__clkbuf_2
Xfanout326 _09564_/A vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__buf_2
Xfanout337 _12441_/S vssd1 vssd1 vccd1 vccd1 _12443_/S sky130_fd_sc_hd__buf_8
X_09813_ _09987_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout348 _08912_/S vssd1 vssd1 vccd1 vccd1 _08932_/S sky130_fd_sc_hd__buf_8
Xfanout359 _15507_/Y vssd1 vssd1 vccd1 vccd1 _15560_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ _09936_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09675_ _10191_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__or2_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _12444_/A hold587/X vssd1 vssd1 vccd1 vccd1 _15935_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _09015_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _15902_/D sky130_fd_sc_hd__and2_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _14774_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_212_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_397_wb_clk_i clkbuf_6_36_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ hold3982/X _10646_/B _10449_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_326_wb_clk_i clkbuf_6_46_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17903_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09109_ hold2102/X _09119_/A2 _09108_/X _12990_/A vssd1 vssd1 vccd1 vccd1 _09109_/X
+ sky130_fd_sc_hd__o211a_1
X_10381_ hold3882/X _10477_/A2 _10380_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _10381_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _12261_/A _12120_/B vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12051_ _12051_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__or2_1
Xhold380 hold380/A vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold391 hold391/A vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ hold4827/X _11192_/B _11001_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout860 _13864_/A vssd1 vssd1 vccd1 vccd1 _13825_/A sky130_fd_sc_hd__buf_8
Xfanout871 fanout873/X vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__buf_8
X_15810_ _17689_/CLK _15810_/D vssd1 vssd1 vccd1 vccd1 _15810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout882 hold1107/X vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__buf_4
X_16790_ _18059_/CLK _16790_/D vssd1 vssd1 vccd1 vccd1 _16790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout893 hold926/X vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__buf_8
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _17712_/CLK _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfxtp_1
X_12953_ hold3253/X _12952_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12954_/B sky130_fd_sc_hd__mux2_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1080 hold1080/A vssd1 vssd1 vccd1 vccd1 _15121_/A sky130_fd_sc_hd__buf_12
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1091 _09306_/X vssd1 vssd1 vccd1 vccd1 _16263_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _13797_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_213_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18460_ _18460_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
X_15672_ _17164_/CLK _15672_/D vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12884_ hold3145/X _12883_/X _12986_/S vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__mux2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ hold1757/X _14612_/B _14622_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14623_/X
+ sky130_fd_sc_hd__o211a_1
X_17411_ _17413_/CLK _17411_/D vssd1 vssd1 vccd1 vccd1 _17411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18391_ _18391_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
X_11835_ _12024_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__or2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17343_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _17342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14554_ hold6005/X _14535_/B hold809/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 hold810/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ hold5068/X _11670_/A _11765_/X vssd1 vssd1 vccd1 vccd1 _11766_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13505_ hold1059/X hold5459/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__mux2_1
X_10717_ hold4403/X _11762_/B _10716_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _10717_/X
+ sky130_fd_sc_hd__o211a_1
X_17273_ _17273_/CLK _17273_/D vssd1 vssd1 vccd1 vccd1 _17273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14485_ _15545_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _11706_/A _11697_/B vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16224_ _18432_/CLK _16224_/D vssd1 vssd1 vccd1 vccd1 _16224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ hold3019/X hold5689/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10648_ _11218_/A _10648_/B vssd1 vssd1 vccd1 vccd1 _16706_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ _17509_/CLK _16155_/D vssd1 vssd1 vccd1 vccd1 _16155_/Q sky130_fd_sc_hd__dfxtp_1
X_13367_ hold2461/X hold3306/X _13847_/C vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__mux2_1
X_10579_ _10603_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _16683_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15106_ hold2755/X _15113_/B _15105_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _15106_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12318_ hold4691/X _12285_/A _12317_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16086_ _18410_/CLK _16086_/D vssd1 vssd1 vccd1 vccd1 hold549/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _17588_/Q _17122_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__mux2_1
X_15037_ _14984_/A hold3092/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12249_ _12273_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__or2_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2709 _17964_/Q vssd1 vssd1 vccd1 vccd1 hold2709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07790_ hold531/X vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__inv_2
X_16988_ _17834_/CLK _16988_/D vssd1 vssd1 vccd1 vccd1 _16988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _17286_/CLK _15939_/D vssd1 vssd1 vccd1 vccd1 hold562/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09460_ _09463_/C _09463_/D _09463_/B vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_235_1382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08411_ _15525_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08411_/X sky130_fd_sc_hd__or2_1
X_17609_ _17641_/CLK _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ hold5856/A _09342_/B _09342_/Y _09390_/X _12404_/A vssd1 vssd1 vccd1 vccd1
+ _09391_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_231_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ hold915/X hold1128/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ hold1515/X _08268_/B _08272_/X _12750_/A vssd1 vssd1 vccd1 vccd1 _08273_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6003 _15835_/Q vssd1 vssd1 vccd1 vccd1 hold6003/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6014 data_in[6] vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6025 _16516_/Q vssd1 vssd1 vccd1 vccd1 hold6025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6036 _16310_/Q vssd1 vssd1 vccd1 vccd1 hold6036/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6047 _16531_/Q vssd1 vssd1 vccd1 vccd1 hold6047/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5302 _16864_/Q vssd1 vssd1 vccd1 vccd1 hold5302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5313 _10297_/X vssd1 vssd1 vccd1 vccd1 _16589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5324 _16614_/Q vssd1 vssd1 vccd1 vccd1 hold5324/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5335 _11545_/X vssd1 vssd1 vccd1 vccd1 _17005_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4601 hold6039/X vssd1 vssd1 vccd1 vccd1 hold4601/X sky130_fd_sc_hd__clkbuf_2
Xhold5346 _17190_/Q vssd1 vssd1 vccd1 vccd1 hold5346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4612 _16349_/Q vssd1 vssd1 vccd1 vccd1 _13262_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5357 _12124_/X vssd1 vssd1 vccd1 vccd1 _17198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4623 _16347_/Q vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5368 _16877_/Q vssd1 vssd1 vccd1 vccd1 hold5368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4634 _16520_/Q vssd1 vssd1 vccd1 vccd1 hold4634/X sky130_fd_sc_hd__buf_2
Xhold5379 _16763_/Q vssd1 vssd1 vccd1 vccd1 hold5379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3900 _16405_/Q vssd1 vssd1 vccd1 vccd1 hold3900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4645 _17100_/Q vssd1 vssd1 vccd1 vccd1 hold4645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4656 _17096_/Q vssd1 vssd1 vccd1 vccd1 hold4656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3911 _11341_/X vssd1 vssd1 vccd1 vccd1 _16937_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3922 _16823_/Q vssd1 vssd1 vccd1 vccd1 hold3922/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4667 _11160_/Y vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4678 hold6038/X vssd1 vssd1 vccd1 vccd1 hold4678/X sky130_fd_sc_hd__buf_1
Xhold3933 _11338_/X vssd1 vssd1 vccd1 vccd1 _16936_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3944 _16595_/Q vssd1 vssd1 vccd1 vccd1 hold3944/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4689 _16923_/Q vssd1 vssd1 vccd1 vccd1 hold4689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3955 _10342_/X vssd1 vssd1 vccd1 vccd1 _16604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3966 _16392_/Q vssd1 vssd1 vccd1 vccd1 hold3966/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3977 _09823_/X vssd1 vssd1 vccd1 vccd1 _16431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout156 _12974_/S vssd1 vssd1 vccd1 vccd1 _12986_/S sky130_fd_sc_hd__buf_4
Xhold3988 _17572_/Q vssd1 vssd1 vccd1 vccd1 hold3988/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout167 _13808_/B vssd1 vssd1 vccd1 vccd1 _13817_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3999 _11533_/X vssd1 vssd1 vccd1 vccd1 _17001_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout178 _11747_/B vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__buf_4
X_07988_ _15557_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
Xfanout189 _12052_/A2 vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__buf_4
XFILLER_0_199_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ hold4006/X _10010_/B _09726_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09658_ hold4819/X _11177_/B _09657_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _09658_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08609_ hold17/X hold235/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_195_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ hold3708/X _10565_/B _09588_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09589_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ hold5184/X _12308_/B _11619_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11620_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ hold5212/X _11747_/B _11550_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ hold1612/X hold4849/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14270_ _15004_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__nand2_1
X_11482_ hold3486/X _11584_/A2 _11481_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11482_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_160_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13221_ _13220_/X hold4655/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__mux2_1
X_10433_ hold3053/X _16635_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _13145_/X _13151_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17537_/D sky130_fd_sc_hd__o21a_1
X_10364_ hold2465/X _16612_/Q _11096_/S vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ hold4913/X _13811_/B _12102_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _12103_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5880 hold5880/A vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_12
X_17960_ _17960_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13082_/X _16903_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10295_ hold3095/X _16589_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__mux2_1
Xhold5891 _18422_/Q vssd1 vssd1 vccd1 vccd1 hold5891/X sky130_fd_sc_hd__dlygate4sd3_1
X_12034_ hold5128/X _13798_/A2 _12033_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12034_/X
+ sky130_fd_sc_hd__o211a_1
X_16911_ _17885_/CLK _16911_/D vssd1 vssd1 vccd1 vccd1 _16911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_236_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17891_ _17891_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16842_ _18430_/CLK _16842_/D vssd1 vssd1 vccd1 vccd1 _16842_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout690 _14442_/C1 vssd1 vssd1 vccd1 vccd1 _14374_/A sky130_fd_sc_hd__buf_4
XFILLER_0_232_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16773_ _18038_/CLK _16773_/D vssd1 vssd1 vccd1 vccd1 _16773_/Q sky130_fd_sc_hd__dfxtp_1
X_13985_ hold2711/X _13986_/B _13984_/Y _13919_/A vssd1 vssd1 vccd1 vccd1 _13985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15724_ _17695_/CLK _15724_/D vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _12999_/A _12936_/B vssd1 vssd1 vccd1 vccd1 _17488_/D sky130_fd_sc_hd__and2_1
XFILLER_0_220_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18443_ _18445_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15655_ _17199_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _12870_/A _12867_/B vssd1 vssd1 vccd1 vccd1 _17465_/D sky130_fd_sc_hd__and2_1
XFILLER_0_197_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _14946_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__nand2_1
X_11818_ hold4976/X _13811_/B _11817_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _11818_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18374_ _18374_/CLK hold857/X vssd1 vssd1 vccd1 vccd1 hold856/A sky130_fd_sc_hd__dfxtp_1
X_15586_ _17200_/CLK _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_248_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18186_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ _12810_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _17442_/D sky130_fd_sc_hd__and2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _18423_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _17325_/Q sky130_fd_sc_hd__dfxtp_1
X_14537_ _14878_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14537_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11749_ _13864_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _17073_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14468_ hold3220/X _14482_/A2 _14467_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17256_ _18447_/CLK _17256_/D vssd1 vssd1 vccd1 vccd1 _17256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13419_ _13713_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13419_/X sky130_fd_sc_hd__or2_1
X_16207_ _18434_/CLK _16207_/D vssd1 vssd1 vccd1 vccd1 _16207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17187_ _17283_/CLK _17187_/D vssd1 vssd1 vccd1 vccd1 _17187_/Q sky130_fd_sc_hd__dfxtp_1
X_14399_ _14794_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _17313_/CLK _16138_/D vssd1 vssd1 vccd1 vccd1 hold544/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _09015_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _16097_/D sky130_fd_sc_hd__and2_1
X_16069_ _17314_/CLK _16069_/D vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__dfxtp_1
Xhold3207 _18381_/Q vssd1 vssd1 vccd1 vccd1 hold3207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3218 _12803_/X vssd1 vssd1 vccd1 vccd1 _12804_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3229 _17450_/Q vssd1 vssd1 vccd1 vccd1 hold3229/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2506 _15719_/Q vssd1 vssd1 vccd1 vccd1 hold2506/X sky130_fd_sc_hd__dlygate4sd3_1
X_07911_ hold2929/X _07918_/B _07910_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07911_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2517 _14777_/X vssd1 vssd1 vccd1 vccd1 _18177_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08891_ _15304_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__and2_1
Xhold2528 _09201_/X vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 _07987_/X vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _18237_/Q vssd1 vssd1 vccd1 vccd1 hold1805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 _09425_/X vssd1 vssd1 vccd1 vccd1 _16298_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07842_ hold1540/X _07865_/B _07841_/X _08119_/A vssd1 vssd1 vccd1 vccd1 _07842_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1827 _18256_/Q vssd1 vssd1 vccd1 vccd1 hold1827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1838 _14396_/X vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 _16318_/Q vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__dlygate4sd3_1
X_09512_ hold940/X _13094_/A _10004_/C vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_211_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09447_/C _09447_/D _09442_/Y vssd1 vssd1 vccd1 vccd1 _09443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ hold477/X _15485_/A2 _15485_/B1 hold674/X _09373_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ _15549_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _14529_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08187_ _14246_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08187_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5110 _16458_/Q vssd1 vssd1 vccd1 vccd1 hold5110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5121 _11302_/X vssd1 vssd1 vccd1 vccd1 _16924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5132 _17257_/Q vssd1 vssd1 vccd1 vccd1 hold5132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5143 _10807_/X vssd1 vssd1 vccd1 vccd1 _16759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5154 _16896_/Q vssd1 vssd1 vccd1 vccd1 hold5154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4420 _10816_/X vssd1 vssd1 vccd1 vccd1 _16762_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5165 _11104_/X vssd1 vssd1 vccd1 vccd1 _16858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_219_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5176 _16472_/Q vssd1 vssd1 vccd1 vccd1 hold5176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4431 _17059_/Q vssd1 vssd1 vccd1 vccd1 hold4431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4442 _13498_/X vssd1 vssd1 vccd1 vccd1 _17619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5187 _11923_/X vssd1 vssd1 vccd1 vccd1 _17131_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5198 _16496_/Q vssd1 vssd1 vccd1 vccd1 hold5198/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4453 _16764_/Q vssd1 vssd1 vccd1 vccd1 hold4453/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4464 _11707_/X vssd1 vssd1 vccd1 vccd1 _17059_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3730 _17430_/Q vssd1 vssd1 vccd1 vccd1 hold3730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4475 _17281_/Q vssd1 vssd1 vccd1 vccd1 hold4475/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3741 _13878_/Y vssd1 vssd1 vccd1 vccd1 _13879_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10080_ _10470_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10080_/X sky130_fd_sc_hd__or2_1
Xhold4486 _11959_/X vssd1 vssd1 vccd1 vccd1 _17143_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3752 _16567_/Q vssd1 vssd1 vccd1 vccd1 hold3752/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4497 _17746_/Q vssd1 vssd1 vccd1 vccd1 hold4497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3763 _11332_/X vssd1 vssd1 vccd1 vccd1 _16934_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_238_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3774 _17159_/Q vssd1 vssd1 vccd1 vccd1 hold3774/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3785 _17408_/Q vssd1 vssd1 vccd1 vccd1 hold3785/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3796 _12671_/X vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13776_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__or2_1
X_10982_ hold2951/X _16818_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12721_ hold2585/X _17418_/Q _12751_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15440_ _15985_/Q _09365_/B _09362_/D _16124_/Q _15438_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_194_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12652_ hold1499/X hold3661/X _12763_/S vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_341_wb_clk_i clkbuf_6_43_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17746_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11603_ hold1763/X hold4319/X _12344_/C vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__mux2_1
X_15371_ _16301_/Q _15477_/A2 _15487_/B1 hold111/X _15370_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/D sky130_fd_sc_hd__a221o_1
X_12583_ hold2614/X _17372_/Q _12967_/S vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14322_ _14878_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__nand2_1
X_17110_ _17270_/CLK _17110_/D vssd1 vssd1 vccd1 vccd1 _17110_/Q sky130_fd_sc_hd__dfxtp_1
X_18090_ _18154_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
X_11534_ hold2068/X _17002_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17041_ _17887_/CLK _17041_/D vssd1 vssd1 vccd1 vccd1 _17041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ hold3165/X _14272_/B _14252_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11465_ hold2258/X hold5581/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ hold4632/X _13203_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__mux2_1
X_10416_ _10536_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14184_ _15203_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14184_/X sky130_fd_sc_hd__or2_1
X_11396_ hold2430/X _16956_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ _13199_/A1 _13133_/X _13134_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13135_/X
+ sky130_fd_sc_hd__o211a_1
X_10347_ _10830_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _17559_/Q _17093_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__mux2_1
X_17943_ _18039_/CLK _17943_/D vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10278_ _10560_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12017_ hold2719/X _17163_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17874_ _17897_/CLK _17874_/D vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
X_16825_ _18058_/CLK _16825_/D vssd1 vssd1 vccd1 vccd1 _16825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756_ _18053_/CLK _16756_/D vssd1 vssd1 vccd1 vccd1 _16756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13968_ _15529_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_429_wb_clk_i clkbuf_6_11_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_216_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _17261_/CLK _15707_/D vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__dfxtp_1
X_12919_ hold1587/X hold3294/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__mux2_1
X_16687_ _18153_/CLK _16687_/D vssd1 vssd1 vccd1 vccd1 _16687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13899_ _14374_/A _13899_/B vssd1 vssd1 vccd1 vccd1 _17755_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_236_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18426_ _18426_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15638_ _17234_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _18389_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15569_ _17274_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _14116_/A hold2534/X hold240/X vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__mux2_1
X_17308_ _17340_/CLK _17308_/D vssd1 vssd1 vccd1 vccd1 hold620/A sky130_fd_sc_hd__dfxtp_1
X_09090_ _15531_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _18350_/CLK hold981/X vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08041_ _14782_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08041_/X sky130_fd_sc_hd__or2_1
X_17239_ _17777_/CLK _17239_/D vssd1 vssd1 vccd1 vccd1 _17239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold902 hold902/A vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold913 hold995/X vssd1 vssd1 vccd1 vccd1 hold996/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 hold935/X vssd1 vssd1 vccd1 vccd1 hold936/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold935 la_data_in[4] vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold946 hold946/A vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3004 _18089_/Q vssd1 vssd1 vccd1 vccd1 hold3004/X sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _16488_/Q _10013_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__and3_1
XFILLER_0_40_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3015 _18282_/Q vssd1 vssd1 vccd1 vccd1 hold3015/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold979 input49/X vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3026 _14811_/X vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ hold88/X hold111/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__mux2_1
Xhold3037 _14478_/X vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3048 _14625_/X vssd1 vssd1 vccd1 vccd1 _18104_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2303 _07925_/X vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3059 _17930_/Q vssd1 vssd1 vccd1 vccd1 hold3059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 _17776_/Q vssd1 vssd1 vccd1 vccd1 hold2314/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2325 _15870_/Q vssd1 vssd1 vccd1 vccd1 hold2325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2336 _07963_/X vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _15021_/X vssd1 vssd1 vccd1 vccd1 _15022_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ hold215/X hold473/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__mux2_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2347 _16221_/Q vssd1 vssd1 vccd1 vccd1 hold2347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1613 _14855_/X vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _08069_/X vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _17804_/Q vssd1 vssd1 vccd1 vccd1 hold1624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _17790_/Q vssd1 vssd1 vccd1 vccd1 hold2369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1635 _14530_/X vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 _18327_/Q vssd1 vssd1 vccd1 vccd1 hold1646/X sky130_fd_sc_hd__dlygate4sd3_1
X_07825_ _07809_/X _07810_/Y hold2013/X _09362_/A vssd1 vssd1 vccd1 vccd1 _07825_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _14029_/X vssd1 vssd1 vccd1 vccd1 _17818_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 _17864_/Q vssd1 vssd1 vccd1 vccd1 hold1668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 _14971_/X vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _09438_/B _16299_/Q vssd1 vssd1 vccd1 vccd1 _09426_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ _09357_/A _09357_/B vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08308_ hold2070/X _08323_/B _08307_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08308_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09288_ hold1618/X _09338_/A2 _09287_/X _12606_/A vssd1 vssd1 vccd1 vccd1 _09288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08239_ hold2199/X _08263_/A2 _08238_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11637_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10201_ hold5316/X _10619_/B _10200_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10201_/X
+ sky130_fd_sc_hd__o211a_1
X_11181_ hold4614/X _11100_/A _11180_/X vssd1 vssd1 vccd1 vccd1 _11181_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4250 _15343_/X vssd1 vssd1 vccd1 vccd1 _15344_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10132_ hold3754/X _10628_/B _10131_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _10132_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4261 _17138_/Q vssd1 vssd1 vccd1 vccd1 hold4261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4272 _15243_/X vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4283 _16807_/Q vssd1 vssd1 vccd1 vccd1 hold4283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4294 _11506_/X vssd1 vssd1 vccd1 vccd1 _16992_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3560 _10011_/Y vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10063_ _10603_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _16511_/D sky130_fd_sc_hd__nor2_1
XTAP_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3571 _16544_/Q vssd1 vssd1 vccd1 vccd1 hold3571/X sky130_fd_sc_hd__dlygate4sd3_1
X_14940_ _15209_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14940_/X sky130_fd_sc_hd__or2_1
XFILLER_0_237_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3582 _10611_/Y vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3593 _17362_/Q vssd1 vssd1 vccd1 vccd1 hold3593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2870 _08420_/X vssd1 vssd1 vccd1 vccd1 _15840_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ hold1773/X _14882_/B _14870_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14871_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2881 _07836_/X vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_214_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2892 _18051_/Q vssd1 vssd1 vccd1 vccd1 hold2892/X sky130_fd_sc_hd__dlygate4sd3_1
X_16610_ _18166_/CLK _16610_/D vssd1 vssd1 vccd1 vccd1 _16610_/Q sky130_fd_sc_hd__dfxtp_1
X_13822_ _13825_/A _13822_/B vssd1 vssd1 vccd1 vccd1 _17727_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_173_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17590_ _17590_/CLK _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16541_ _18181_/CLK _16541_/D vssd1 vssd1 vccd1 vccd1 _16541_/Q sky130_fd_sc_hd__dfxtp_1
X_13753_ hold4533/X _13847_/B _13752_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ _11061_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ hold3779/X _12703_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16472_ _18383_/CLK _16472_/D vssd1 vssd1 vccd1 vccd1 _16472_/Q sky130_fd_sc_hd__dfxtp_1
X_13684_ hold4259/X _13886_/B _13683_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10896_ _11094_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18211_ _18231_/CLK hold875/X vssd1 vssd1 vccd1 vccd1 hold874/A sky130_fd_sc_hd__dfxtp_1
X_15423_ _15481_/A1 _15415_/X _15422_/X _15481_/B1 hold5874/A vssd1 vssd1 vccd1 vccd1
+ _15423_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ hold3336/X _12634_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ _15394_/A _15354_/B vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__and2_1
X_18142_ _18142_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ hold3472/X _12565_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14305_ hold3073/X hold756/X _14304_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11517_ _12285_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ _15285_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15285_/X sky130_fd_sc_hd__or2_1
X_18073_ _18108_/CLK hold916/X vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
X_12497_ hold14/X _12509_/A2 _12507_/A3 _12496_/X _09053_/A vssd1 vssd1 vccd1 vccd1
+ hold15/A sky130_fd_sc_hd__o311a_1
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 input23/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__buf_1
X_14236_ _15185_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17024_ _17905_/CLK _17024_/D vssd1 vssd1 vccd1 vccd1 _17024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11448_ _11553_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ hold1545/X _14198_/B _14166_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _11667_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__or2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _15551_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14098_/X sky130_fd_sc_hd__or2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold5859/X hold960/X _13055_/C vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17926_ _17960_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17889_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_240_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16808_ _18041_/CLK _16808_/D vssd1 vssd1 vccd1 vccd1 _16808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08590_ hold292/X hold828/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold829/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_263_wb_clk_i clkbuf_6_56_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17968_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17788_ _17883_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ _18068_/CLK _16739_/D vssd1 vssd1 vccd1 vccd1 _16739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09211_ hold2748/X _09216_/B _09210_/X _12894_/A vssd1 vssd1 vccd1 vccd1 _09211_/X
+ sky130_fd_sc_hd__o211a_1
X_18409_ _18409_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09142_ _15525_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ hold1176/X _09119_/A2 _09072_/X _12999_/A vssd1 vssd1 vccd1 vccd1 _09073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08024_ hold2800/X _08029_/B _08023_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08024_/X
+ sky130_fd_sc_hd__o211a_1
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold721 hold721/A vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold732 hold732/A vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold754 hold754/A vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold765 hold765/A vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__buf_2
Xhold776 hold776/A vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 hold787/A vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _10467_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__or2_1
Xhold798 hold798/A vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2100 _15728_/Q vssd1 vssd1 vccd1 vccd1 hold2100/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2111 _14569_/X vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ hold140/X hold356/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__mux2_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2122 _14571_/X vssd1 vssd1 vccd1 vccd1 _18078_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _14173_/X vssd1 vssd1 vccd1 vccd1 _17887_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2144 _12970_/X vssd1 vssd1 vccd1 vccd1 hold2144/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _15663_/Q vssd1 vssd1 vccd1 vccd1 hold1410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 _17762_/Q vssd1 vssd1 vccd1 vccd1 hold2155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2166 _15578_/Q vssd1 vssd1 vccd1 vccd1 hold2166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 _14005_/X vssd1 vssd1 vccd1 vccd1 _17806_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08857_ _12418_/A hold218/X vssd1 vssd1 vccd1 vccd1 _16047_/D sky130_fd_sc_hd__and2_1
XFILLER_0_157_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2177 _14771_/X vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 _18431_/Q vssd1 vssd1 vccd1 vccd1 hold1432/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1443 _14237_/X vssd1 vssd1 vccd1 vccd1 _17917_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2188 _18447_/Q vssd1 vssd1 vccd1 vccd1 hold2188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2199 _15754_/Q vssd1 vssd1 vccd1 vccd1 hold2199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 _17784_/Q vssd1 vssd1 vccd1 vccd1 hold1454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1465 _09127_/X vssd1 vssd1 vccd1 vccd1 _16176_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07808_ _12412_/A _13048_/A _07803_/Y hold2045/X vssd1 vssd1 vccd1 vccd1 _07808_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1476 _17975_/Q vssd1 vssd1 vccd1 vccd1 hold1476/X sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ _15454_/A hold317/X vssd1 vssd1 vccd1 vccd1 _16014_/D sky130_fd_sc_hd__and2_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _15853_/Q vssd1 vssd1 vccd1 vccd1 hold1487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _14991_/X vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10750_ hold5477/X _11732_/B _10749_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10750_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09409_ _07804_/A _09447_/B _15264_/A _09408_/X vssd1 vssd1 vccd1 vccd1 _09409_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ hold5415/X _11159_/B _10680_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _10681_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12420_ _12424_/A hold831/X vssd1 vssd1 vccd1 vccd1 _17303_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ hold3602/X _13461_/A _12350_/X vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_wb_clk_i clkbuf_6_25_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18460_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11302_ hold5120/X _12314_/B _11301_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__o211a_1
X_15070_ _15070_/A hold623/X vssd1 vssd1 vccd1 vccd1 hold624/A sky130_fd_sc_hd__and2_1
XFILLER_0_205_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _13782_/A _12282_/B vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__or2_1
XFILLER_0_239_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ hold993/X _14040_/B _14020_/X _15500_/A vssd1 vssd1 vccd1 vccd1 hold994/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ hold3831/X _11617_/A2 _11232_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11164_ _11203_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _16878_/D sky130_fd_sc_hd__nor2_1
XTAP_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4080 _11824_/X vssd1 vssd1 vccd1 vccd1 _17098_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_234_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ hold2397/X hold4725/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4091 _17162_/Q vssd1 vssd1 vccd1 vccd1 hold4091/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _17299_/CLK _15972_/D vssd1 vssd1 vccd1 vccd1 hold813/A sky130_fd_sc_hd__dfxtp_1
X_11095_ _11189_/A _11095_/A2 _11094_/X _14667_/C1 vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ _17711_/CLK _17711_/D vssd1 vssd1 vccd1 vccd1 _17711_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3390 _17480_/Q vssd1 vssd1 vccd1 vccd1 hold3390/X sky130_fd_sc_hd__dlygate4sd3_1
X_14923_ hold6001/X _14946_/B hold927/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 hold928/A
+ sky130_fd_sc_hd__o211a_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _16506_/Q _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__and3_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17642_ _17642_/CLK _17642_/D vssd1 vssd1 vccd1 vccd1 _17642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _14854_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _17722_/Q _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13805_/X sky130_fd_sc_hd__and3_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ _17739_/CLK _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
X_14785_ hold1555/X _14772_/B _14784_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14785_/X
+ sky130_fd_sc_hd__o211a_1
X_11997_ _13794_/A _11997_/B vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ _18176_/CLK _16524_/D vssd1 vssd1 vccd1 vccd1 _16524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_1406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ hold3444/X _11729_/B _10947_/X _14554_/C1 vssd1 vssd1 vccd1 vccd1 _10948_/X
+ sky130_fd_sc_hd__o211a_1
X_13736_ hold2100/X hold5727/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16455_ _18366_/CLK _16455_/D vssd1 vssd1 vccd1 vccd1 _16455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10879_ hold5050/X _11168_/B _10878_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__o211a_1
X_13667_ hold1662/X _17676_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15406_ _17344_/Q _15448_/B1 _15485_/B1 hold92/X vssd1 vssd1 vccd1 vccd1 _15406_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _12870_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _17382_/D sky130_fd_sc_hd__and2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _18391_/CLK _16386_/D vssd1 vssd1 vccd1 vccd1 _16386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13598_ hold1474/X hold3462/X _13874_/C vssd1 vssd1 vccd1 vccd1 _13599_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _18213_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15337_ hold489/X _15487_/A2 _15484_/B1 hold506/X _15336_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/B sky130_fd_sc_hd__a221o_2
X_12549_ _13002_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _17359_/D sky130_fd_sc_hd__and2_1
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5709 _17694_/Q vssd1 vssd1 vccd1 vccd1 hold5709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_26_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_26_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_18056_ _18065_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _13057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ hold617/X _09386_/A _15451_/A2 hold629/X vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17007_ _17885_/CLK _17007_/D vssd1 vssd1 vccd1 vccd1 _17007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ hold1939/X _14216_/Y _14218_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15199_ _15199_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout508 _10400_/S vssd1 vssd1 vccd1 vccd1 _10565_/C sky130_fd_sc_hd__clkbuf_8
Xfanout519 _09499_/Y vssd1 vssd1 vccd1 vccd1 _10025_/C sky130_fd_sc_hd__buf_12
XFILLER_0_10_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09760_ hold4851/X _10049_/B _09759_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_225_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_444_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08711_ hold263/X hold460/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold461/A sky130_fd_sc_hd__mux2_1
XFILLER_0_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17909_ _18070_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09691_ hold4723/X _10601_/B _09690_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08642_ _15264_/A hold229/X vssd1 vssd1 vccd1 vccd1 _15943_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08573_ _12416_/A hold354/X vssd1 vssd1 vccd1 vccd1 _15910_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09125_ _15128_/A hold533/X vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__or2_2
XFILLER_0_162_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09056_ hold140/X _16145_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08007_ _15521_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08007_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 data_in[0] vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold562 hold562/A vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold573/A vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 hold584/A vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 input34/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09958_ _10052_/A _10468_/A2 _09957_/X _15226_/C1 vssd1 vssd1 vccd1 vccd1 _09958_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_185_wb_clk_i clkbuf_6_54_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18108_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _12426_/A hold849/X vssd1 vssd1 vccd1 vccd1 _16072_/D sky130_fd_sc_hd__and2_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_6_21_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17523_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09889_ hold3370/X _10025_/B _09888_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1240 _07874_/X vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 _08255_/X vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ hold4091/X _13811_/B _11919_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _11920_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1262 _15512_/X vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_213_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1273 _18253_/Q vssd1 vssd1 vccd1 vccd1 hold1273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 _14983_/X vssd1 vssd1 vccd1 vccd1 _18275_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1295 _07967_/X vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ hold5306/X _12347_/B _11850_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ hold2190/X hold5086/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__mux2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14570_ hold690/X _14573_/B hold2120/X vssd1 vssd1 vccd1 vccd1 _14570_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _13864_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _17084_/D sky130_fd_sc_hd__nor2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ hold2512/X _16735_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13521_ _13713_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13452_ _13761_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__or2_1
X_16240_ _18445_/CLK _16240_/D vssd1 vssd1 vccd1 vccd1 _16240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ hold1038/X hold3679/X _11156_/C vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ hold361/X hold868/X _12441_/S vssd1 vssd1 vccd1 vccd1 hold869/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _13794_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_1
X_16171_ _17508_/CLK _16171_/D vssd1 vssd1 vccd1 vccd1 _16171_/Q sky130_fd_sc_hd__dfxtp_1
X_10595_ _16689_/Q _10619_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15122_ hold1232/X _15113_/B _15121_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _15122_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ _13873_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _17268_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ hold469/X hold471/X _15071_/S vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__mux2_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ hold4115/X _13868_/B _12264_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12265_/X
+ sky130_fd_sc_hd__o211a_1
X_14004_ hold915/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__or2_1
X_11216_ _16896_/Q _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__and3_1
XFILLER_0_31_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12196_ hold5234/X _13798_/A2 _12195_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput82 _13209_/A vssd1 vssd1 vccd1 vccd1 output82/X sky130_fd_sc_hd__buf_6
Xoutput93 _13289_/A vssd1 vssd1 vccd1 vccd1 output93/X sky130_fd_sc_hd__buf_6
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11147_ _16873_/Q _11147_/B _11147_/C vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__and3_1
XFILLER_0_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15955_ _17322_/CLK _15955_/D vssd1 vssd1 vccd1 vccd1 hold413/A sky130_fd_sc_hd__dfxtp_1
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ hold2892/X _16850_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_223_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10029_ _13190_/A _09954_/A _10028_/X vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__a21oi_1
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ hold926/X _14910_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or2_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _17160_/CLK _15886_/D vssd1 vssd1 vccd1 vccd1 _15886_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17625_ _17689_/CLK _17625_/D vssd1 vssd1 vccd1 vccd1 _17625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14837_ hold1229/X _14828_/B _14836_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14837_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _18221_/CLK _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14768_ _14946_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ _18322_/CLK _16507_/D vssd1 vssd1 vccd1 vccd1 _16507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _13800_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13719_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17487_ _17508_/CLK _17487_/D vssd1 vssd1 vccd1 vccd1 _17487_/Q sky130_fd_sc_hd__dfxtp_1
X_14699_ hold3141/X _14714_/B _14698_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16438_ _18349_/CLK _16438_/D vssd1 vssd1 vccd1 vccd1 _16438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16369_ _18376_/CLK _16369_/D vssd1 vssd1 vccd1 vccd1 _16369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18108_ _18108_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5506 _11392_/X vssd1 vssd1 vccd1 vccd1 _16954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5517 _16786_/Q vssd1 vssd1 vccd1 vccd1 hold5517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5528 _09928_/X vssd1 vssd1 vccd1 vccd1 _16466_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5539 _16798_/Q vssd1 vssd1 vccd1 vccd1 hold5539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4805 _16611_/Q vssd1 vssd1 vccd1 vccd1 hold4805/X sky130_fd_sc_hd__dlygate4sd3_1
X_18039_ _18039_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4816 _11763_/Y vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4827 _16856_/Q vssd1 vssd1 vccd1 vccd1 hold4827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4838 _09742_/X vssd1 vssd1 vccd1 vccd1 _16404_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4849 _16658_/Q vssd1 vssd1 vccd1 vccd1 hold4849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout305 _09984_/A vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__buf_4
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout316 _11094_/A vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__buf_4
Xfanout327 _10476_/A vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__buf_4
X_09812_ hold1102/X _16428_/Q _10004_/C vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__mux2_1
Xfanout338 _12401_/S vssd1 vssd1 vccd1 vccd1 _12441_/S sky130_fd_sc_hd__buf_8
XFILLER_0_22_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout349 _08793_/S vssd1 vssd1 vccd1 vccd1 _08779_/S sky130_fd_sc_hd__buf_8
XFILLER_0_226_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09743_ hold2479/X _16405_/Q _10007_/C vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ hold2927/X hold5669/X _10190_/S vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ hold454/X hold586/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold587/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ hold271/X hold342/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08487_ hold1735/X _08486_/B _08486_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 _08487_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _15549_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10380_ _10476_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ _12436_/A hold476/X vssd1 vssd1 vccd1 vccd1 _16136_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_366_wb_clk_i clkbuf_6_34_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17647_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ hold2282/X hold5473/X _12338_/C vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold381 hold381/A vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 hold392/A vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__buf_4
X_11001_ _11097_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout850 _15215_/A vssd1 vssd1 vccd1 vccd1 _14946_/A sky130_fd_sc_hd__buf_12
Xfanout861 _13864_/A vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__buf_8
XFILLER_0_217_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout872 fanout873/X vssd1 vssd1 vccd1 vccd1 _18461_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout883 hold1107/X vssd1 vssd1 vccd1 vccd1 hold1108/A sky130_fd_sc_hd__clkbuf_1
Xfanout894 hold925/X vssd1 vssd1 vccd1 vccd1 hold926/A sky130_fd_sc_hd__buf_6
X_15740_ _17744_/CLK _15740_/D vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ hold968/X hold3244/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__mux2_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 _18248_/Q vssd1 vssd1 vccd1 vccd1 hold1070/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _15067_/X vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 _18383_/Q vssd1 vssd1 vccd1 vccd1 hold1092/X sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ hold1243/X hold5134/X _13412_/S vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15671_ _17195_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ hold2806/X _17472_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux2_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17431_/CLK _17410_/D vssd1 vssd1 vccd1 vccd1 _17410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _15231_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14622_/X sky130_fd_sc_hd__or2_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18390_/CLK hold888/X vssd1 vssd1 vccd1 vccd1 hold887/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11834_ hold2534/X hold4653/X _13862_/C vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17341_ _17346_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _17341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14553_ hold808/X _14553_/B vssd1 vssd1 vccd1 vccd1 hold809/A sky130_fd_sc_hd__or2_1
X_11765_ _17079_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_6_16_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17496_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _11667_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__or2_1
X_13504_ hold3462/X _13880_/B _13503_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13504_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17272_ _17272_/CLK _17272_/D vssd1 vssd1 vccd1 vccd1 _17272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_6_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17258_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11696_ hold2624/X _17056_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__mux2_1
X_14484_ hold2075/X _14487_/B _14483_/Y _14554_/C1 vssd1 vssd1 vccd1 vccd1 _14484_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ _17455_/CLK _16223_/D vssd1 vssd1 vccd1 vccd1 _16223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10647_ hold3607/X _10998_/A _10646_/X vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__a21oi_1
X_13435_ hold4934/X _13817_/B _13434_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ _17491_/CLK _16154_/D vssd1 vssd1 vccd1 vccd1 _16154_/Q sky130_fd_sc_hd__dfxtp_1
X_13366_ hold4269/X _12374_/B _13365_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _13366_/X
+ sky130_fd_sc_hd__o211a_1
X_10578_ hold4601/X _10482_/A _10577_/X vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ _15105_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15105_/X sky130_fd_sc_hd__or2_1
X_12317_ _17263_/Q _12317_/B _12317_/C vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__and3_1
X_13297_ _13297_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13297_/X sky130_fd_sc_hd__and2_1
X_16085_ _18407_/CLK _16085_/D vssd1 vssd1 vccd1 vccd1 hold639/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15036_ _15058_/A _15036_/B vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__and2_1
X_12248_ hold2286/X _17240_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12179_ hold2667/X _17217_/Q _13556_/S vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16987_ _17842_/CLK _16987_/D vssd1 vssd1 vccd1 vccd1 _16987_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _17301_/CLK _15938_/D vssd1 vssd1 vccd1 vccd1 hold410/A sky130_fd_sc_hd__dfxtp_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15869_ _17612_/CLK _15869_/D vssd1 vssd1 vccd1 vccd1 _15869_/Q sky130_fd_sc_hd__dfxtp_1
X_08410_ hold6003/X _08440_/A2 hold1010/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_235_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ _17738_/CLK _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_1
X_09390_ _09369_/C _09389_/X _18458_/Q vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _08391_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _15802_/D sky130_fd_sc_hd__and2_1
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17539_ _18378_/CLK _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08272_ _15551_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08272_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6004 _16319_/Q vssd1 vssd1 vccd1 vccd1 hold6004/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6015 _18417_/Q vssd1 vssd1 vccd1 vccd1 hold6015/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6026 _17522_/Q vssd1 vssd1 vccd1 vccd1 hold960/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6037 _15854_/Q vssd1 vssd1 vccd1 vccd1 hold6037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5303 _11026_/X vssd1 vssd1 vccd1 vccd1 _16832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6048 _16308_/Q vssd1 vssd1 vccd1 vccd1 hold6048/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5314 _17007_/Q vssd1 vssd1 vccd1 vccd1 hold5314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5325 _10276_/X vssd1 vssd1 vccd1 vccd1 _16582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5336 _16780_/Q vssd1 vssd1 vccd1 vccd1 hold5336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4602 _16346_/Q vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5347 _12004_/X vssd1 vssd1 vccd1 vccd1 _17158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4613 _10056_/Y vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5358 _17135_/Q vssd1 vssd1 vccd1 vccd1 hold5358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4624 _10050_/Y vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5369 _11065_/X vssd1 vssd1 vccd1 vccd1 _16845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4635 _10569_/Y vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3901 _09649_/X vssd1 vssd1 vccd1 vccd1 _16373_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4646 _12309_/Y vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4657 _12297_/Y vssd1 vssd1 vccd1 vccd1 _12298_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3912 _17001_/Q vssd1 vssd1 vccd1 vccd1 hold3912/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4668 _16354_/Q vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3923 _10903_/X vssd1 vssd1 vccd1 vccd1 _16791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3934 _16944_/Q vssd1 vssd1 vccd1 vccd1 hold3934/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4679 _16904_/Q vssd1 vssd1 vccd1 vccd1 hold4679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3945 _10219_/X vssd1 vssd1 vccd1 vccd1 _16563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3956 _16641_/Q vssd1 vssd1 vccd1 vccd1 hold3956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3967 _09610_/X vssd1 vssd1 vccd1 vccd1 _16360_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3978 _17274_/Q vssd1 vssd1 vccd1 vccd1 hold3978/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout157 _12965_/S vssd1 vssd1 vccd1 vccd1 _13001_/S sky130_fd_sc_hd__buf_6
Xhold3989 _13836_/Y vssd1 vssd1 vccd1 vccd1 _13837_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout168 _12031_/A2 vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__clkbuf_8
X_07987_ hold2538/X _07978_/B _07986_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _07987_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout179 _11150_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09726_ _09933_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__or2_1
XFILLER_0_215_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09657_ _11082_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _12416_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _15926_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _10560_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__or2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _09055_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _15893_/D sky130_fd_sc_hd__and2_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ _12285_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11550_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ hold5425/X _10619_/B _10500_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11481_ _11679_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ hold4625/X _13219_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__mux2_1
X_10432_ hold3787/X _10622_/B _10431_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151_ _13199_/A1 _13149_/X _13150_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13151_/X
+ sky130_fd_sc_hd__o211a_1
X_10363_ hold4978/X _10649_/B _10362_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12102_ _13716_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__or2_1
X_13082_ _17561_/Q _17095_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__mux2_1
Xhold5870 hold5870/A vssd1 vssd1 vccd1 vccd1 hold5870/X sky130_fd_sc_hd__clkbuf_4
Xhold5881 _18418_/Q vssd1 vssd1 vccd1 vccd1 hold5881/X sky130_fd_sc_hd__dlygate4sd3_1
X_10294_ hold3908/X _10622_/B _10293_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5892 hold5892/A vssd1 vssd1 vccd1 vccd1 hold5892/X sky130_fd_sc_hd__clkbuf_4
X_12033_ _12288_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__or2_1
X_16910_ _17852_/CLK _16910_/D vssd1 vssd1 vccd1 vccd1 _16910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17890_ _17890_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _18042_/CLK _16841_/D vssd1 vssd1 vccd1 vccd1 _16841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_232_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout680 _15494_/A vssd1 vssd1 vccd1 vccd1 _14149_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_219_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout691 fanout692/X vssd1 vssd1 vccd1 vccd1 _14442_/C1 sky130_fd_sc_hd__clkbuf_4
X_16772_ _18071_/CLK _16772_/D vssd1 vssd1 vccd1 vccd1 _16772_/Q sky130_fd_sc_hd__dfxtp_1
X_13984_ _15545_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15723_ _17157_/CLK _15723_/D vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ hold3269/X _12934_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12936_/B sky130_fd_sc_hd__mux2_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18442_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15654_ _17198_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12866_ hold3325/X _12865_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__mux2_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ hold2955/X _14612_/B _14604_/X _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14605_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18373_ _18373_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ _13716_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__or2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _17164_/CLK _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ hold3337/X _12796_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__mux2_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _18411_/CLK hold27/X vssd1 vssd1 vccd1 vccd1 _17324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ hold2323/X _14535_/B _14535_/Y _13921_/A vssd1 vssd1 vccd1 vccd1 _14536_/X
+ sky130_fd_sc_hd__o211a_1
X_11748_ hold3583/X _12219_/A _11747_/X vssd1 vssd1 vccd1 vccd1 _11748_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _17444_/CLK _17255_/D vssd1 vssd1 vccd1 vccd1 _17255_/Q sky130_fd_sc_hd__dfxtp_1
X_14467_ _15201_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11679_ _11679_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_288_wb_clk_i clkbuf_6_37_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18050_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ _18434_/CLK _16206_/D vssd1 vssd1 vccd1 vccd1 _16206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13418_ hold2715/X hold3424/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17186_ _17639_/CLK _17186_/D vssd1 vssd1 vccd1 vccd1 _17186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14398_ hold1393/X _14446_/A2 _14397_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _14398_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_217_wb_clk_i clkbuf_6_60_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18205_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16137_ _17332_/CLK _16137_/D vssd1 vssd1 vccd1 vccd1 hold428/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ hold1138/X hold5657/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3208 _15202_/X vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16068_ _17299_/CLK _16068_/D vssd1 vssd1 vccd1 vccd1 hold852/A sky130_fd_sc_hd__dfxtp_1
Xhold3219 _17503_/Q vssd1 vssd1 vccd1 vccd1 hold3219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ hold2927/X hold514/X _15018_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15019_/X
+ sky130_fd_sc_hd__o211a_1
X_07910_ _15533_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__or2_1
Xhold2507 _18300_/Q vssd1 vssd1 vccd1 vccd1 hold2507/X sky130_fd_sc_hd__dlygate4sd3_1
X_08890_ hold98/X hold847/X _08928_/S vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__mux2_1
Xhold2518 _18449_/Q vssd1 vssd1 vccd1 vccd1 hold2518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2529 _17824_/Q vssd1 vssd1 vccd1 vccd1 hold2529/X sky130_fd_sc_hd__dlygate4sd3_1
X_07841_ _14854_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__or2_1
XFILLER_0_237_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1806 _14903_/X vssd1 vssd1 vccd1 vccd1 _18237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1817 _16314_/Q vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_236_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1828 _14943_/X vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 _18196_/Q vssd1 vssd1 vccd1 vccd1 hold1839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09511_ hold3384/X _10013_/B _09510_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _09511_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09442_ _09447_/C _09447_/D _09484_/B vssd1 vssd1 vccd1 vccd1 _09442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09373_ _17325_/Q _15487_/A2 _15487_/B1 hold678/X vssd1 vssd1 vccd1 vccd1 _09373_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08324_ hold2085/X _08336_/A2 _08323_/Y _08367_/A vssd1 vssd1 vccd1 vccd1 _08324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ hold5977/X _08263_/A2 hold1250/X _08389_/A vssd1 vssd1 vccd1 vccd1 _08255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08186_ hold1567/X _08209_/B _08185_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5100 _17164_/Q vssd1 vssd1 vccd1 vccd1 hold5100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5111 _09808_/X vssd1 vssd1 vccd1 vccd1 _16426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5122 _16934_/Q vssd1 vssd1 vccd1 vccd1 hold5122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5133 _12205_/X vssd1 vssd1 vccd1 vccd1 _17225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5144 _16849_/Q vssd1 vssd1 vccd1 vccd1 hold5144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5155 _11122_/X vssd1 vssd1 vccd1 vccd1 _16864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4410 _11863_/X vssd1 vssd1 vccd1 vccd1 _17111_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5166 _16854_/Q vssd1 vssd1 vccd1 vccd1 hold5166/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4421 _16990_/Q vssd1 vssd1 vccd1 vccd1 hold4421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5177 _09850_/X vssd1 vssd1 vccd1 vccd1 _16440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4432 _11611_/X vssd1 vssd1 vccd1 vccd1 _17027_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4443 _17027_/Q vssd1 vssd1 vccd1 vccd1 hold4443/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5188 _16790_/Q vssd1 vssd1 vccd1 vccd1 hold5188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5199 _09922_/X vssd1 vssd1 vccd1 vccd1 _16464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4454 _10726_/X vssd1 vssd1 vccd1 vccd1 _16732_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4465 _17606_/Q vssd1 vssd1 vccd1 vccd1 hold4465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3720 _16732_/Q vssd1 vssd1 vccd1 vccd1 hold3720/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3731 _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4476 _12277_/X vssd1 vssd1 vccd1 vccd1 _17249_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3742 _16592_/Q vssd1 vssd1 vccd1 vccd1 hold3742/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4487 _16977_/Q vssd1 vssd1 vccd1 vccd1 hold4487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3753 _10135_/X vssd1 vssd1 vccd1 vccd1 _16535_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4498 _13783_/X vssd1 vssd1 vccd1 vccd1 _17714_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3764 _16624_/Q vssd1 vssd1 vccd1 vccd1 hold3764/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3775 _11911_/X vssd1 vssd1 vccd1 vccd1 _17127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_233_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3786 _17412_/Q vssd1 vssd1 vccd1 vccd1 hold3786/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3797 _16655_/Q vssd1 vssd1 vccd1 vccd1 hold3797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ hold3357/X _10013_/B _09708_/X _15186_/C1 vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10981_ hold5144/X _11738_/B _10980_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _10981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _12759_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _17416_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ _12654_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _17393_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11602_ hold4437/X _11801_/B _11601_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15370_ hold676/X _15486_/A2 _09357_/B _16066_/Q vssd1 vssd1 vccd1 vccd1 _15370_/X
+ sky130_fd_sc_hd__a22o_1
X_12582_ _12969_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _17370_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ hold2583/X _14326_/B _14320_/Y _14667_/C1 vssd1 vssd1 vccd1 vccd1 _14321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ hold3998/X _11726_/B _11532_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11533_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_381_wb_clk_i clkbuf_6_33_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17040_ _17886_/CLK _17040_/D vssd1 vssd1 vccd1 vccd1 _17040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _15201_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__or2_1
X_11464_ hold5338/X _11738_/B _11463_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11464_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_310_wb_clk_i clkbuf_6_45_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17994_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_208_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10415_ hold1935/X hold3793/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__mux2_1
X_13203_ _13202_/X _16918_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ hold5326/X _12317_/B _11394_/X _14013_/C1 vssd1 vssd1 vccd1 vccd1 _11395_/X
+ sky130_fd_sc_hd__o211a_1
X_14183_ hold2683/X _14202_/B _14182_/X _14472_/C1 vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ _13134_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__or2_1
X_10346_ hold2812/X hold3920/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__and2_1
X_17942_ _18045_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ hold3141/X hold4835/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12016_ hold4917/X _12293_/B _12015_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _12016_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17873_ _17905_/CLK _17873_/D vssd1 vssd1 vccd1 vccd1 _17873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16824_ _18200_/CLK _16824_/D vssd1 vssd1 vccd1 vccd1 _16824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16755_ _18319_/CLK _16755_/D vssd1 vssd1 vccd1 vccd1 _16755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ hold3057/X _13995_/A2 _13966_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_221_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15706_ _17178_/CLK _15706_/D vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _12921_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _17482_/D sky130_fd_sc_hd__and2_1
X_16686_ _18210_/CLK _16686_/D vssd1 vssd1 vccd1 vccd1 _16686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13898_ _15513_/A hold2642/X hold124/X vssd1 vssd1 vccd1 vccd1 _13899_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18425_ _18425_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15637_ _17266_/CLK _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12849_ _12870_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _17459_/D sky130_fd_sc_hd__and2_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18356_ _18356_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15568_ _17639_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ _17327_/CLK _17307_/D vssd1 vssd1 vccd1 vccd1 _17307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14519_ _14984_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18287_ _18287_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
X_15499_ _15515_/A hold1972/X hold691/X vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08040_ hold2486/X _08033_/B _08039_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _08040_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17238_ _17767_/CLK _17238_/D vssd1 vssd1 vccd1 vccd1 _17238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 hold997/X vssd1 vssd1 vccd1 vccd1 hold998/A sky130_fd_sc_hd__buf_6
X_17169_ _17266_/CLK _17169_/D vssd1 vssd1 vccd1 vccd1 _17169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold925 hold937/X vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 hold936/A vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 la_data_in[9] vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _11203_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _16487_/D sky130_fd_sc_hd__nor2_1
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3005 _14595_/X vssd1 vssd1 vccd1 vccd1 _18089_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3016 _14997_/X vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3027 _18186_/Q vssd1 vssd1 vccd1 vccd1 hold3027/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3038 _18308_/Q vssd1 vssd1 vccd1 vccd1 hold3038/X sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ _15364_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _16088_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2304 _16155_/Q vssd1 vssd1 vccd1 vccd1 hold2304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3049 _16210_/Q vssd1 vssd1 vccd1 vccd1 hold3049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _15792_/Q vssd1 vssd1 vccd1 vccd1 hold2315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _08483_/X vssd1 vssd1 vccd1 vccd1 _15870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2337 _17783_/Q vssd1 vssd1 vccd1 vccd1 hold2337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ _12416_/A hold420/X vssd1 vssd1 vccd1 vccd1 _16054_/D sky130_fd_sc_hd__and2_1
Xhold1603 _16275_/Q vssd1 vssd1 vccd1 vccd1 hold1603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _09219_/X vssd1 vssd1 vccd1 vccd1 _16221_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1614 _16189_/Q vssd1 vssd1 vccd1 vccd1 hold1614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2359 _15744_/Q vssd1 vssd1 vccd1 vccd1 hold2359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1625 _13999_/X vssd1 vssd1 vccd1 vccd1 _17804_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07824_ _09366_/A _09122_/A _07824_/C _09121_/B vssd1 vssd1 vccd1 vccd1 _07824_/Y
+ sky130_fd_sc_hd__nor4_2
Xhold1636 _17929_/Q vssd1 vssd1 vccd1 vccd1 hold1636/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1647 _15090_/X vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1658 _17918_/Q vssd1 vssd1 vccd1 vccd1 hold1658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1669 _14125_/X vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ _07785_/Y hold5972/X _15304_/A _09424_/X vssd1 vssd1 vccd1 vccd1 _09425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_220_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _09366_/A _09366_/B _09356_/C vssd1 vssd1 vccd1 vccd1 _09356_/Y sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_139_wb_clk_i clkbuf_6_31_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17534_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _15531_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09287_ _14968_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08238_ _14403_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08169_ _15500_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _10524_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ _16884_/Q _11180_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__and3_1
XTAP_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4240 _16825_/Q vssd1 vssd1 vccd1 vccd1 hold4240/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ _10497_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__or2_1
Xhold4251 _17652_/Q vssd1 vssd1 vccd1 vccd1 hold4251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4262 _11848_/X vssd1 vssd1 vccd1 vccd1 _17106_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4273 _17282_/Q vssd1 vssd1 vccd1 vccd1 hold4273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4284 _10855_/X vssd1 vssd1 vccd1 vccd1 _16775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3550 _10614_/Y vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4295 _16754_/Q vssd1 vssd1 vccd1 vccd1 hold4295/X sky130_fd_sc_hd__dlygate4sd3_1
X_10062_ _13278_/A _10488_/A _10061_/X vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_234_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3561 _17378_/Q vssd1 vssd1 vccd1 vccd1 hold3561/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3572 _10641_/Y vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3583 _16913_/Q vssd1 vssd1 vccd1 vccd1 hold3583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3594 _12557_/X vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2860 _17880_/Q vssd1 vssd1 vccd1 vccd1 hold2860/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2871 _18297_/Q vssd1 vssd1 vccd1 vccd1 hold2871/X sky130_fd_sc_hd__dlygate4sd3_1
X_14870_ _15209_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__or2_1
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2882 _16216_/Q vssd1 vssd1 vccd1 vccd1 hold2882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 _14514_/X vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13821_ hold5659/X _13734_/A _13820_/X vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _18212_/CLK _16540_/D vssd1 vssd1 vccd1 vccd1 _16540_/Q sky130_fd_sc_hd__dfxtp_1
X_13752_ _13776_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__or2_1
X_10964_ hold2705/X _16812_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ hold2179/X _17412_/Q _12763_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _18382_/CLK _16471_/D vssd1 vssd1 vccd1 vccd1 _16471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13683_ _13779_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10895_ hold2664/X _16789_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18210_ _18210_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15422_ _15480_/A _15422_/B _15422_/C _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_156_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12634_ hold1237/X hold3331/X _12772_/S vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _18141_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
X_15353_ _15481_/A1 _15345_/X _15352_/X _15481_/B1 _18409_/Q vssd1 vssd1 vccd1 vccd1
+ _15353_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_136_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12565_ hold3002/X _17366_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14304_ _14984_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14304_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18072_ _18078_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11516_ hold2409/X hold3930/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15284_ _15324_/A _15284_/B vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__and2_1
Xclkbuf_6_16_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_16_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _17341_/Q _12498_/B vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17023_ _17869_/CLK _17023_/D vssd1 vssd1 vccd1 vccd1 _17023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ hold1593/X _14266_/B _14234_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14235_/X
+ sky130_fd_sc_hd__o211a_1
X_11447_ hold2821/X _16973_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14166_ hold915/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14166_/X sky130_fd_sc_hd__or2_1
X_11378_ hold2058/X _16950_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13117_ _13116_/X hold4601/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_10329_ _10830_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__or2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ hold2271/X _14094_/B _14096_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14097_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13048_ _13048_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__and2_1
X_17925_ _18063_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ _17888_/CLK _17856_/D vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16807_ _18040_/CLK _16807_/D vssd1 vssd1 vccd1 vccd1 _16807_/Q sky130_fd_sc_hd__dfxtp_1
X_17787_ _17851_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
X_14999_ hold1398/X hold514/X _14998_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ _17971_/CLK _16738_/D vssd1 vssd1 vccd1 vccd1 _16738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16669_ _18225_/CLK _16669_/D vssd1 vssd1 vccd1 vccd1 _16669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_6_55_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_55_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09210_ _15539_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__or2_1
X_18408_ _18408_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_232_wb_clk_i clkbuf_6_63_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18219_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ hold1423/X _09177_/A2 _09140_/X _12912_/A vssd1 vssd1 vccd1 vccd1 _09141_/X
+ sky130_fd_sc_hd__o211a_1
X_18339_ _18397_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09072_ _14972_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08023_ _15537_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08023_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold700 hold700/A vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 hold711/A vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold722 hold722/A vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold733 hold733/A vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__clkbuf_8
Xhold744 hold744/A vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold755 hold755/A vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__buf_2
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/A vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 hold788/A vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ hold1470/X hold5094/X _10190_/S vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2101 _08184_/X vssd1 vssd1 vccd1 vccd1 _15728_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2112 _17972_/Q vssd1 vssd1 vccd1 vccd1 hold2112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2123 hold2140/X vssd1 vssd1 vccd1 vccd1 hold2141/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08925_ _15414_/A hold157/X vssd1 vssd1 vccd1 vccd1 _16080_/D sky130_fd_sc_hd__and2_1
XFILLER_0_239_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2134 _18451_/Q vssd1 vssd1 vccd1 vccd1 hold2134/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_239_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2145 _12971_/X vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 la_data_in[10] vssd1 vssd1 vccd1 vccd1 hold1400/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2156 _15645_/Q vssd1 vssd1 vccd1 vccd1 hold2156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 _08044_/X vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1422 _16228_/Q vssd1 vssd1 vccd1 vccd1 hold1422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 _07866_/X vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ hold210/X hold217/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__mux2_1
Xhold1433 _15510_/X vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2178 _16248_/Q vssd1 vssd1 vccd1 vccd1 hold2178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2189 _15542_/X vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 _15562_/Q vssd1 vssd1 vccd1 vccd1 hold1444/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1455 _13959_/X vssd1 vssd1 vccd1 vccd1 _17784_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 _18358_/Q vssd1 vssd1 vccd1 vccd1 hold1466/X sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ _07785_/Y _07789_/A _07805_/A _07806_/Y vssd1 vssd1 vccd1 vccd1 _07807_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1477 _15690_/Q vssd1 vssd1 vccd1 vccd1 hold1477/X sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ hold140/X hold316/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__mux2_1
Xhold1488 _08446_/X vssd1 vssd1 vccd1 vccd1 _15853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _18444_/Q vssd1 vssd1 vccd1 vccd1 hold1499/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09408_ _09438_/B _16290_/Q vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__or2_1
X_10680_ _11064_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09339_ _09339_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_36_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _17274_/Q _12374_/B _13556_/S vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__and3_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _12219_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12281_ hold2560/X hold4289/X _13877_/C vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14020_ hold944/X _14042_/B vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__or2_1
X_11232_ _11712_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ hold4699/X _11106_/A _11162_/X vssd1 vssd1 vccd1 vccd1 _11163_/Y sky130_fd_sc_hd__a21oi_1
XTAP_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_6_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17816_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4070 _11251_/X vssd1 vssd1 vccd1 vccd1 _16907_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ hold3748/X _10628_/B _10113_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10114_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4081 _17597_/Q vssd1 vssd1 vccd1 vccd1 hold4081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ _18408_/CLK _15971_/D vssd1 vssd1 vccd1 vccd1 hold789/A sky130_fd_sc_hd__dfxtp_1
X_11094_ _11094_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4092 _11920_/X vssd1 vssd1 vccd1 vccd1 _17130_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3380 _09919_/X vssd1 vssd1 vccd1 vccd1 _16463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17710_ _17742_/CLK _17710_/D vssd1 vssd1 vccd1 vccd1 _17710_/Q sky130_fd_sc_hd__dfxtp_1
X_10045_ _10603_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _16505_/D sky130_fd_sc_hd__nor2_1
XTAP_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ hold926/X _14964_/B vssd1 vssd1 vccd1 vccd1 hold927/A sky130_fd_sc_hd__or2_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3391 _17479_/Q vssd1 vssd1 vccd1 vccd1 hold3391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__clkbuf_1
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2690 _14695_/X vssd1 vssd1 vccd1 vccd1 _18137_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _17641_/CLK _17641_/D vssd1 vssd1 vccd1 vccd1 _17641_/Q sky130_fd_sc_hd__dfxtp_1
X_14853_ hold2443/X _14880_/B _14852_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14853_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_215_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13825_/A _13804_/B vssd1 vssd1 vccd1 vccd1 _17721_/D sky130_fd_sc_hd__nor2_1
X_17572_ _17680_/CLK _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
X_14784_ _15231_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14784_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11996_ hold1542/X hold4158/X _12029_/S vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__mux2_1
X_16523_ _18143_/CLK _16523_/D vssd1 vssd1 vccd1 vccd1 _16523_/Q sky130_fd_sc_hd__dfxtp_1
X_13735_ hold5705/X _13829_/B _13734_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _11637_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__or2_1
XFILLER_0_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ _18397_/CLK _16454_/D vssd1 vssd1 vccd1 vccd1 _16454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13666_ hold4376/X _13856_/B _13665_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13666_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _11553_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10878_/X sky130_fd_sc_hd__or2_1
X_15405_ hold609/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12617_ hold3415/X _12616_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_213_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16385_ _16517_/CLK _16385_/D vssd1 vssd1 vccd1 vccd1 _16385_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ hold4255/X _13883_/B _13596_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13597_/X
+ sky130_fd_sc_hd__o211a_1
X_18124_ _18124_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
X_15336_ _17337_/Q _15448_/B1 _15485_/B1 hold516/X vssd1 vssd1 vccd1 vccd1 _15336_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ hold3588/X _12547_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18055_ _18055_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ hold632/X _15487_/A2 _09386_/D hold322/X _15266_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/B sky130_fd_sc_hd__a221o_1
X_12479_ hold35/X _12445_/A _12445_/B _12478_/X _12438_/A vssd1 vssd1 vccd1 vccd1
+ hold36/A sky130_fd_sc_hd__o311a_1
XANTENNA_2 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17006_ _17884_/CLK _17006_/D vssd1 vssd1 vccd1 vccd1 _17006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ _14968_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14218_/X sky130_fd_sc_hd__or2_1
X_15198_ hold1481/X _15221_/B _15197_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _15198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_238_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ hold2278/X _14148_/B _14148_/Y _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14149_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout509 _10481_/S vssd1 vssd1 vccd1 vccd1 _10055_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08710_ _12404_/A hold900/X vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__and2_1
X_17908_ _17908_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09690_ _10488_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__or2_1
XFILLER_0_222_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08641_ hold228/X _15943_/Q _08655_/S vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__mux2_1
XFILLER_0_238_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _17871_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_234_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ hold353/X _15910_/Q _08594_/S vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_413_wb_clk_i clkbuf_6_14_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17897_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ _15128_/A hold533/X vssd1 vssd1 vccd1 vccd1 _09124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_199_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09055_/A hold425/X vssd1 vssd1 vccd1 vccd1 _16144_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08006_ hold1542/X _08029_/B _08005_/X _08115_/A vssd1 vssd1 vccd1 vccd1 _08006_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold530 input60/X vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold552 hold79/X vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 hold563/A vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold574 hold574/A vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 hold71/X vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__buf_4
XFILLER_0_217_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _10191_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__or2_1
XFILLER_0_217_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ hold402/X hold848/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold849/A sky130_fd_sc_hd__mux2_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _09984_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__or2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _14837_/X vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _15686_/Q vssd1 vssd1 vccd1 vccd1 hold1241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 _16170_/Q vssd1 vssd1 vccd1 vccd1 hold1252/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _15304_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _16038_/D sky130_fd_sc_hd__and2_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1263 _18021_/Q vssd1 vssd1 vccd1 vccd1 hold1263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _14937_/X vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _15652_/Q vssd1 vssd1 vccd1 vccd1 hold1285/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _16276_/Q vssd1 vssd1 vccd1 vccd1 hold1296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _12231_/A _11850_/B vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_154_wb_clk_i clkbuf_6_28_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ hold5168/X _11216_/B _10800_/X _14542_/C1 vssd1 vssd1 vccd1 vccd1 _10801_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ hold4662/X _12219_/A _11780_/X vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ hold2596/X hold4032/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ hold5549/X _11762_/B _10731_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10732_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ hold1652/X _17604_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10663_ hold4407/X _11147_/B _10662_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10663_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12402_ _15324_/A hold671/X vssd1 vssd1 vccd1 vccd1 _17294_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _17507_/CLK _16170_/D vssd1 vssd1 vccd1 vccd1 _16170_/Q sky130_fd_sc_hd__dfxtp_1
X_10594_ _11194_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _16688_/D sky130_fd_sc_hd__nor2_1
X_13382_ hold2325/X hold4747/X _13793_/S vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__mux2_1
X_15121_ _15121_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12333_ hold3611/X _13773_/A _12332_/X vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15052_ _15052_/A _15052_/B vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12264_ _13773_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14003_ hold1704/X _14038_/B _14002_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14003_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11215_ _11218_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _16895_/D sky130_fd_sc_hd__nor2_1
X_12195_ _13797_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput72 _13051_/A vssd1 vssd1 vccd1 vccd1 output72/X sky130_fd_sc_hd__buf_6
Xoutput83 _13065_/A vssd1 vssd1 vccd1 vccd1 output83/X sky130_fd_sc_hd__buf_6
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11146_ _11158_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _16872_/D sky130_fd_sc_hd__nor2_1
Xoutput94 _13073_/A vssd1 vssd1 vccd1 vccd1 output94/X sky130_fd_sc_hd__buf_6
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15954_ _17286_/CLK _15954_/D vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__dfxtp_1
X_11077_ hold5084/X _11738_/B _11076_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _11077_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10028_ _10028_/A _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__and3_1
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _18238_/Q _14896_/Y hold1336/X _15482_/A vssd1 vssd1 vccd1 vccd1 _14905_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _17723_/CLK _15885_/D vssd1 vssd1 vccd1 vccd1 _15885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _15121_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14836_/X sky130_fd_sc_hd__or2_1
X_17624_ _17694_/CLK _17624_/D vssd1 vssd1 vccd1 vccd1 _17624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17555_ _18131_/CLK _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14767_ hold1921/X _14774_/B _14766_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14767_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _12267_/A _11979_/B vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16506_ _18360_/CLK _16506_/D vssd1 vssd1 vccd1 vccd1 _16506_/Q sky130_fd_sc_hd__dfxtp_1
X_13718_ hold1622/X hold3395/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17486_ _17508_/CLK _17486_/D vssd1 vssd1 vccd1 vccd1 _17486_/Q sky130_fd_sc_hd__dfxtp_1
X_14698_ _14984_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16437_ _18316_/CLK _16437_/D vssd1 vssd1 vccd1 vccd1 _16437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13649_ hold1096/X _17670_/Q _13841_/C vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16368_ _18377_/CLK _16368_/D vssd1 vssd1 vccd1 vccd1 _16368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _18263_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_1
X_15319_ _15973_/Q _15485_/A2 _15488_/A2 hold434/X _15318_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5507 _17022_/Q vssd1 vssd1 vccd1 vccd1 hold5507/X sky130_fd_sc_hd__dlygate4sd3_1
X_16299_ _16320_/CLK _16299_/D vssd1 vssd1 vccd1 vccd1 _16299_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5518 _10792_/X vssd1 vssd1 vccd1 vccd1 _16754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5529 _17043_/Q vssd1 vssd1 vccd1 vccd1 hold5529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _18038_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4806 _10267_/X vssd1 vssd1 vccd1 vccd1 _16579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4817 _16507_/Q vssd1 vssd1 vccd1 vccd1 hold4817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4828 _11002_/X vssd1 vssd1 vccd1 vccd1 _16824_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4839 _16634_/Q vssd1 vssd1 vccd1 vccd1 hold4839/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout306 _11061_/A vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__buf_4
X_09811_ hold4034/X _10007_/B _09810_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09811_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout317 fanout334/X vssd1 vssd1 vccd1 vccd1 _11094_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout328 _10476_/A vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout339 _09369_/X vssd1 vssd1 vccd1 vccd1 _15483_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ hold4837/X _10049_/B _09741_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09742_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ hold4767/X _10055_/B _09672_/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 _09673_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _15414_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _15934_/D sky130_fd_sc_hd__and2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _12424_/A hold802/X vssd1 vssd1 vccd1 vccd1 _15901_/D sky130_fd_sc_hd__and2_1
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08486_ _15004_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ hold2184/X _09106_/B _09106_/Y _12987_/A vssd1 vssd1 vccd1 vccd1 _09107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ hold402/X hold475/X _09056_/S vssd1 vssd1 vccd1 vccd1 hold476/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 input7/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 hold371/A vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold382 hold382/A vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__buf_4
XFILLER_0_229_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold393 hold393/A vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__clkbuf_8
X_11000_ hold2721/X hold4781/X _11192_/C vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout840 fanout847/X vssd1 vssd1 vccd1 vccd1 _14839_/C1 sky130_fd_sc_hd__buf_4
Xfanout851 _07783_/Y vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__buf_12
Xfanout862 fanout873/X vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__buf_8
Xfanout873 input71/X vssd1 vssd1 vccd1 vccd1 fanout873/X sky130_fd_sc_hd__buf_12
Xfanout884 _15195_/A vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_335_wb_clk_i clkbuf_6_41_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17237_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout895 _14974_/A vssd1 vssd1 vccd1 vccd1 _15515_/A sky130_fd_sc_hd__clkbuf_16
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _12990_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _17493_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _08350_/X vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 _14927_/X vssd1 vssd1 vccd1 vccd1 _18248_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ hold4158/X _12031_/A2 _11901_/X _08155_/A vssd1 vssd1 vccd1 vccd1 _11902_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _15068_/X vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ _17161_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _15206_/X vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _12990_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _17470_/D sky130_fd_sc_hd__and2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ hold2371/X _14612_/B _14620_/X _14797_/C1 vssd1 vssd1 vccd1 vccd1 _14621_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ hold5397/X _13862_/B _11832_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _17340_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 _17340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ hold1960/X _14535_/B _14551_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _12340_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _17078_/D sky130_fd_sc_hd__nor2_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _13791_/A _13503_/B vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__or2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10715_ hold3059/X _16729_/Q _11204_/C vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__mux2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17777_/CLK _17271_/D vssd1 vssd1 vccd1 vccd1 _17271_/Q sky130_fd_sc_hd__dfxtp_1
X_14483_ _15543_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_166_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11695_ hold5613/X _11768_/B _11694_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _11695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16222_ _17455_/CLK _16222_/D vssd1 vssd1 vccd1 vccd1 _16222_/Q sky130_fd_sc_hd__dfxtp_1
X_13434_ _13698_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _13434_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _16706_/Q _10646_/B _10997_/S vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _17491_/CLK _16153_/D vssd1 vssd1 vccd1 vccd1 _16153_/Q sky130_fd_sc_hd__dfxtp_1
X_13365_ _13461_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__or2_1
X_10577_ _10577_/A _10577_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10577_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_6_13_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17882_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15104_ hold2979/X _15113_/B _15103_/X _15192_/C1 vssd1 vssd1 vccd1 vccd1 _15104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _13825_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _17262_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_239_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16084_ _18406_/CLK _16084_/D vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ _13289_/X _13295_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15035_ _15197_/A hold1460/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__mux2_1
X_12247_ hold4529/X _12365_/B _12246_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__o211a_1
X_12178_ hold4370/X _12274_/A2 _12177_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _12178_/X
+ sky130_fd_sc_hd__o211a_1
X_11129_ hold2693/X hold5286/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11130_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _17896_/CLK _16986_/D vssd1 vssd1 vccd1 vccd1 _16986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _17284_/CLK _15937_/D vssd1 vssd1 vccd1 vccd1 hold588/A sky130_fd_sc_hd__dfxtp_1
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _17647_/CLK _15868_/D vssd1 vssd1 vccd1 vccd1 _15868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14819_ hold1937/X _14828_/B _14818_/X _14386_/A vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__o211a_1
X_17607_ _17607_/CLK _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15799_ _17425_/CLK _15799_/D vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08340_ _14164_/A hold1379/X hold134/X vssd1 vssd1 vccd1 vccd1 _08340_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _18378_/CLK _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ hold2214/X _08268_/B _08270_/X _12741_/A vssd1 vssd1 vccd1 vccd1 _08271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17469_ _17469_/CLK _17469_/D vssd1 vssd1 vccd1 vccd1 _17469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6005 _18071_/Q vssd1 vssd1 vccd1 vccd1 hold6005/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6016 _18407_/Q vssd1 vssd1 vccd1 vccd1 hold6016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6027 _17524_/Q vssd1 vssd1 vccd1 vccd1 hold6027/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6038 _16725_/Q vssd1 vssd1 vccd1 vccd1 hold6038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6049 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold6049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5304 _16819_/Q vssd1 vssd1 vccd1 vccd1 hold5304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5315 _11455_/X vssd1 vssd1 vccd1 vccd1 _16975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5326 _16987_/Q vssd1 vssd1 vccd1 vccd1 hold5326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5337 _10774_/X vssd1 vssd1 vccd1 vccd1 _16748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4603 _10047_/Y vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5348 _17165_/Q vssd1 vssd1 vccd1 vccd1 hold5348/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4614 _16724_/Q vssd1 vssd1 vccd1 vccd1 hold4614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5359 _11839_/X vssd1 vssd1 vccd1 vccd1 _17103_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4625 _16728_/Q vssd1 vssd1 vccd1 vccd1 hold4625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4636 hold6047/X vssd1 vssd1 vccd1 vccd1 hold4636/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3902 _16572_/Q vssd1 vssd1 vccd1 vccd1 hold3902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4647 _17564_/Q vssd1 vssd1 vccd1 vccd1 hold4647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4658 _17099_/Q vssd1 vssd1 vccd1 vccd1 hold4658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3913 _11437_/X vssd1 vssd1 vccd1 vccd1 _16969_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4669 _10071_/Y vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3924 _16938_/Q vssd1 vssd1 vccd1 vccd1 hold3924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3935 _11266_/X vssd1 vssd1 vccd1 vccd1 _16912_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3946 _16428_/Q vssd1 vssd1 vccd1 vccd1 hold3946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3957 _10357_/X vssd1 vssd1 vccd1 vccd1 _16609_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3968 _16358_/Q vssd1 vssd1 vccd1 vccd1 hold3968/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout147 _12755_/S vssd1 vssd1 vccd1 vccd1 _12764_/S sky130_fd_sc_hd__buf_6
Xfanout158 _12968_/S vssd1 vssd1 vccd1 vccd1 _12965_/S sky130_fd_sc_hd__buf_6
Xhold3979 _12256_/X vssd1 vssd1 vccd1 vccd1 _17242_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07986_ _15555_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07986_/X sky130_fd_sc_hd__or2_1
Xfanout169 _12031_/A2 vssd1 vssd1 vccd1 vccd1 _13862_/B sky130_fd_sc_hd__buf_4
XFILLER_0_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ hold471/X hold3392/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_226_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09656_ hold1043/X _16376_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _09657_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08607_ hold88/X hold93/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__mux2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09587_ hold2685/X _16353_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ hold113/X hold494/X _08592_/S vssd1 vssd1 vccd1 vccd1 _08539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_194_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08469_ hold2195/X _08486_/B _08468_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08469_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10500_ _10524_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ hold2802/X _16984_/Q _11480_/S vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10527_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13150_ _13150_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ _10554_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12101_ hold2640/X hold3837/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5860 hold5860/A vssd1 vssd1 vccd1 vccd1 load_status[5] sky130_fd_sc_hd__buf_12
X_13081_ _13081_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__and2_1
Xhold5871 _18414_/Q vssd1 vssd1 vccd1 vccd1 hold5871/X sky130_fd_sc_hd__dlygate4sd3_1
X_10293_ _10497_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5882 hold5882/A vssd1 vssd1 vccd1 vccd1 hold5882/X sky130_fd_sc_hd__clkbuf_4
Xhold5893 _18415_/Q vssd1 vssd1 vccd1 vccd1 hold5893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ hold2017/X _17168_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__mux2_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16840_ _18041_/CLK _16840_/D vssd1 vssd1 vccd1 vccd1 _16840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout670 _08159_/A vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__buf_4
Xfanout681 _15494_/A vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__buf_4
XFILLER_0_233_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16771_ _18064_/CLK _16771_/D vssd1 vssd1 vccd1 vccd1 _16771_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout692 fanout693/X vssd1 vssd1 vccd1 vccd1 fanout692/X sky130_fd_sc_hd__clkbuf_4
X_13983_ hold2058/X _13986_/B _13982_/Y _13941_/A vssd1 vssd1 vccd1 vccd1 _13983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_219_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15722_ _17129_/CLK _15722_/D vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ hold2568/X hold3267/X _12997_/S vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__mux2_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18441_ _18442_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
X_15653_ _17198_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ hold2096/X hold3303/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__mux2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _15105_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14604_/X sky130_fd_sc_hd__or2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18380_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
X_11816_ hold2019/X hold4656/X _13811_/C vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _17897_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ hold991/X hold3302/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux2_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17323_ _17347_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _17323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14946_/A _14535_/B vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__nand2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _17073_/Q _11747_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17254_ _17254_/CLK _17254_/D vssd1 vssd1 vccd1 vccd1 _17254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14466_ hold3132/X _14487_/B _14465_/X _15194_/C1 vssd1 vssd1 vccd1 vccd1 _14466_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ hold1616/X _17050_/Q _12344_/C vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16205_ _18436_/CLK _16205_/D vssd1 vssd1 vccd1 vccd1 _16205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13417_ hold4101/X _13814_/B _13416_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13417_/X
+ sky130_fd_sc_hd__o211a_1
X_10629_ hold3551/X _10497_/A _10628_/X vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__a21oi_1
X_17185_ _17217_/CLK _17185_/D vssd1 vssd1 vccd1 vccd1 _17185_/Q sky130_fd_sc_hd__dfxtp_1
X_14397_ hold915/X _14411_/B vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16136_ _17335_/CLK _16136_/D vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ hold5753/X _13832_/B _13347_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13348_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _16087_/CLK _16067_/D vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__dfxtp_1
X_13279_ _13311_/A1 _13277_/X _13278_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3209 _17426_/Q vssd1 vssd1 vccd1 vccd1 hold3209/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_257_wb_clk_i clkbuf_6_58_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18054_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15018_ _15233_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2508 _17873_/Q vssd1 vssd1 vccd1 vccd1 hold2508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 _15546_/X vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07840_ hold2182/X _07865_/B _07839_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _07840_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1807 _18455_/Q vssd1 vssd1 vccd1 vccd1 hold1807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1818 _09421_/X vssd1 vssd1 vccd1 vccd1 _16296_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1829 _18190_/Q vssd1 vssd1 vccd1 vccd1 hold1829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16969_ _17815_/CLK _16969_/D vssd1 vssd1 vccd1 vccd1 _16969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09510_ _09918_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__or2_1
XFILLER_0_223_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09441_ _09447_/D _09484_/B vssd1 vssd1 vccd1 vccd1 _16306_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_176_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09372_ _07805_/A _09362_/A _09386_/A hold482/X vssd1 vssd1 vccd1 vccd1 _09375_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ _15547_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _15207_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08185_ _14854_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5101 _11926_/X vssd1 vssd1 vccd1 vccd1 _17132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5112 _16886_/Q vssd1 vssd1 vccd1 vccd1 hold5112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5123 _11236_/X vssd1 vssd1 vccd1 vccd1 _16902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5134 _17125_/Q vssd1 vssd1 vccd1 vccd1 hold5134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5145 _10981_/X vssd1 vssd1 vccd1 vccd1 _16817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4400 _11314_/X vssd1 vssd1 vccd1 vccd1 _16928_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4411 _17283_/Q vssd1 vssd1 vccd1 vccd1 hold4411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5156 _17193_/Q vssd1 vssd1 vccd1 vccd1 hold5156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5167 _10996_/X vssd1 vssd1 vccd1 vccd1 _16822_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4422 _11404_/X vssd1 vssd1 vccd1 vccd1 _16958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5178 _16781_/Q vssd1 vssd1 vccd1 vccd1 hold5178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4433 _17082_/Q vssd1 vssd1 vccd1 vccd1 hold4433/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5189 _10804_/X vssd1 vssd1 vccd1 vccd1 _16758_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4444 _11515_/X vssd1 vssd1 vccd1 vccd1 _16995_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3710 _16683_/Q vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4455 _17674_/Q vssd1 vssd1 vccd1 vccd1 hold4455/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4466 _13363_/X vssd1 vssd1 vccd1 vccd1 _17574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3721 _11205_/Y vssd1 vssd1 vccd1 vccd1 _11206_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3732 _16711_/Q vssd1 vssd1 vccd1 vccd1 hold3732/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4477 _17183_/Q vssd1 vssd1 vccd1 vccd1 hold4477/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3743 _10210_/X vssd1 vssd1 vccd1 vccd1 _16560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4488 _11365_/X vssd1 vssd1 vccd1 vccd1 _16945_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3754 _16566_/Q vssd1 vssd1 vccd1 vccd1 hold3754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4499 _17679_/Q vssd1 vssd1 vccd1 vccd1 hold4499/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3765 _10306_/X vssd1 vssd1 vccd1 vccd1 _16592_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3776 _16675_/Q vssd1 vssd1 vccd1 vccd1 hold3776/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3787 _16666_/Q vssd1 vssd1 vccd1 vccd1 hold3787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3798 _10399_/X vssd1 vssd1 vccd1 vccd1 _16623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ hold2640/X _07978_/B _07968_/X _15548_/C1 vssd1 vssd1 vccd1 vccd1 _07969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_241_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09708_ _09918_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__or2_1
XFILLER_0_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10980_ _11643_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__or2_1
X_09639_ _11106_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ hold3468/X _12649_/X _12755_/S vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_1287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _11706_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12581_ hold3159/X _12580_/X _12968_/S vssd1 vssd1 vccd1 vccd1 _12581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _14946_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ _11631_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ hold3128/X _14266_/B _14250_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11463_ _11643_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _17576_/Q _17110_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__mux2_1
X_10414_ hold4885/X _10649_/B _10413_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14182_ _15201_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14182_/X sky130_fd_sc_hd__or2_1
X_11394_ _12285_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ _13132_/X hold4627/X _13181_/S vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ hold5000/X _10631_/B _10344_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_350_wb_clk_i clkbuf_6_40_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17745_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5690 _13342_/X vssd1 vssd1 vccd1 vccd1 _17567_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13051_/X _13063_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17526_/D sky130_fd_sc_hd__o21a_1
X_17941_ _18014_/CLK hold603/X vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10276_ hold5324/X _10598_/B _10275_/X _14829_/C1 vssd1 vssd1 vccd1 vccd1 _10276_/X
+ sky130_fd_sc_hd__o211a_1
X_12015_ _12288_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17872_ _17872_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16823_ _18230_/CLK _16823_/D vssd1 vssd1 vccd1 vccd1 _16823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_232_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ _15201_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13966_/X sky130_fd_sc_hd__or2_1
X_16754_ _18019_/CLK _16754_/D vssd1 vssd1 vccd1 vccd1 _16754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ _17273_/CLK _15705_/D vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfxtp_1
X_12917_ hold3315/X _12916_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__mux2_1
X_16685_ _18143_/CLK _16685_/D vssd1 vssd1 vccd1 vccd1 _16685_/Q sky130_fd_sc_hd__dfxtp_1
X_13897_ _14376_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _17754_/D sky130_fd_sc_hd__and2_1
XFILLER_0_213_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_6_45_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_45_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_18424_ _18426_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15636_ _17200_/CLK _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ hold3419/X _12847_/X _12914_/S vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18355_ _18379_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15567_ _17895_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ hold3348/X _12778_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17306_ _17306_/CLK _17306_/D vssd1 vssd1 vccd1 vccd1 hold860/A sky130_fd_sc_hd__dfxtp_1
X_14518_ hold1450/X _14541_/B _14517_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18286_ _18390_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14449_ _14968_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__or2_1
X_17237_ _17237_/CLK _17237_/D vssd1 vssd1 vccd1 vccd1 _17237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_438_wb_clk_i clkbuf_6_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17694_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 hold904/A vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _17200_/CLK _17168_/D vssd1 vssd1 vccd1 vccd1 _17168_/Q sky130_fd_sc_hd__dfxtp_1
Xhold915 hold915/A vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__buf_12
Xhold926 hold926/A vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__clkbuf_16
X_16119_ _17343_/CLK _16119_/D vssd1 vssd1 vccd1 vccd1 _16119_/Q sky130_fd_sc_hd__dfxtp_1
Xhold937 input63/X vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 hold948/A vssd1 vssd1 vccd1 vccd1 input68/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _13086_/A _09918_/A _09989_/X vssd1 vssd1 vccd1 vccd1 _09990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17099_ _17195_/CLK _17099_/D vssd1 vssd1 vccd1 vccd1 _17099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3006 _18143_/Q vssd1 vssd1 vccd1 vccd1 hold3006/X sky130_fd_sc_hd__dlygate4sd3_1
X_08941_ hold113/X hold518/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__mux2_1
Xhold3017 _15758_/Q vssd1 vssd1 vccd1 vccd1 hold3017/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3028 _14797_/X vssd1 vssd1 vccd1 vccd1 _18186_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3039 _16184_/Q vssd1 vssd1 vccd1 vccd1 hold3039/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2305 _09081_/X vssd1 vssd1 vccd1 vccd1 _16155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 _08318_/X vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08872_ hold312/X hold419/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold420/A sky130_fd_sc_hd__mux2_1
Xhold2327 _15837_/Q vssd1 vssd1 vccd1 vccd1 hold2327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2338 _13957_/X vssd1 vssd1 vccd1 vccd1 _17783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _09330_/X vssd1 vssd1 vccd1 vccd1 _16275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 _18066_/Q vssd1 vssd1 vccd1 vccd1 hold2349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1615 _09153_/X vssd1 vssd1 vccd1 vccd1 _16189_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07823_ hold246/X hold469/X _09496_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09121_/B
+ sky130_fd_sc_hd__or4b_1
Xhold1626 _17893_/Q vssd1 vssd1 vccd1 vccd1 hold1626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1637 _14261_/X vssd1 vssd1 vccd1 vccd1 _17929_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _18382_/Q vssd1 vssd1 vccd1 vccd1 hold1648/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1659 _14239_/X vssd1 vssd1 vccd1 vccd1 _17918_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ _09438_/B _09424_/B vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _15547_/A _15219_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09356_/C sky130_fd_sc_hd__or3_1
XFILLER_0_136_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08306_ hold1474/X _08336_/A2 _08305_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _08306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09286_ _14913_/A hold533/A vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__or2_2
XFILLER_0_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08237_ hold2445/X _08263_/A2 _08236_/X _13657_/C1 vssd1 vssd1 vccd1 vccd1 _08237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_wb_clk_i clkbuf_6_49_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18387_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08168_ _15519_/A hold1115/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_108_wb_clk_i clkbuf_6_20_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16081_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08099_ hold1186/X _08088_/B _08098_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _08099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4230 _12136_/X vssd1 vssd1 vccd1 vccd1 _17202_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10130_ hold2484/X hold3581/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__mux2_1
Xhold4241 _10909_/X vssd1 vssd1 vccd1 vccd1 _16793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4252 _13501_/X vssd1 vssd1 vccd1 vccd1 _17620_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4263 _17177_/Q vssd1 vssd1 vccd1 vccd1 hold4263/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4274 _12280_/X vssd1 vssd1 vccd1 vccd1 _17250_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3540 _10062_/Y vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4285 _17642_/Q vssd1 vssd1 vccd1 vccd1 hold4285/X sky130_fd_sc_hd__dlygate4sd3_1
X_10061_ _16511_/Q _10577_/B _10481_/S vssd1 vssd1 vccd1 vccd1 _10061_/X sky130_fd_sc_hd__and3_1
XTAP_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3551 _16540_/Q vssd1 vssd1 vccd1 vccd1 hold3551/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4296 _10696_/X vssd1 vssd1 vccd1 vccd1 _16722_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3562 _12605_/X vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3573 _16332_/Q vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3584 _11748_/Y vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2850 _18136_/Q vssd1 vssd1 vccd1 vccd1 hold2850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3595 _17361_/Q vssd1 vssd1 vccd1 vccd1 hold3595/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2861 _14157_/X vssd1 vssd1 vccd1 vccd1 _17880_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2872 _15575_/Q vssd1 vssd1 vccd1 vccd1 hold2872/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2883 _09209_/X vssd1 vssd1 vccd1 vccd1 _16216_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13820_ _17727_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13820_/X sky130_fd_sc_hd__and3_1
Xhold2894 _16164_/Q vssd1 vssd1 vccd1 vccd1 hold2894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ hold2223/X hold4393/X _13841_/C vssd1 vssd1 vccd1 vccd1 _13752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_230_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ hold5485/X _11156_/B _10962_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12702_ _12768_/A _12702_/B vssd1 vssd1 vccd1 vccd1 _17410_/D sky130_fd_sc_hd__and2_1
X_16470_ _18381_/CLK _16470_/D vssd1 vssd1 vccd1 vccd1 _16470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13682_ _15762_/Q _17681_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ hold4785/X _11177_/B _10893_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10894_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ hold792/X _15451_/A2 _09386_/D hold706/X _15416_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_195_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ _12780_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _17387_/D sky130_fd_sc_hd__and2_1
XFILLER_0_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18140_ _18263_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
X_15352_ _15480_/A _15352_/B _15352_/C _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__or4_1
X_12564_ _12960_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _17364_/D sky130_fd_sc_hd__and2_1
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ hold1365/X hold756/X _14302_/X _14370_/A vssd1 vssd1 vccd1 vccd1 _14303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18071_ _18071_/CLK hold810/X vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
X_11515_ hold4443/X _12365_/B _11514_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11515_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15283_ _15490_/A1 _15275_/X _15282_/X _15490_/B1 _18402_/Q vssd1 vssd1 vccd1 vccd1
+ _15283_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_163_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12495_ hold59/X _12445_/A _12445_/B _12494_/X _12430_/A vssd1 vssd1 vccd1 vccd1
+ hold60/A sky130_fd_sc_hd__o311a_1
XFILLER_0_83_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17022_ _17900_/CLK _17022_/D vssd1 vssd1 vccd1 vccd1 _17022_/Q sky130_fd_sc_hd__dfxtp_1
X_14234_ _14968_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ hold4275/X _11729_/B _11445_/X _15496_/A vssd1 vssd1 vccd1 vccd1 _11446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14165_ hold1472/X _14198_/B _14164_/X _14374_/A vssd1 vssd1 vccd1 vccd1 _14165_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ hold5561/X _11768_/B _11376_/X _13921_/A vssd1 vssd1 vccd1 vccd1 _11377_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ hold4903/X _13115_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__mux2_2
X_10328_ hold2878/X hold5082/X _11198_/C vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__mux2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _15549_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13056_/C _13044_/X _13046_/X _09339_/A vssd1 vssd1 vccd1 vccd1 _13047_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17924_ _18319_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ hold1912/X _16577_/Q _10997_/S vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_218_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _17855_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ _18039_/CLK _16806_/D vssd1 vssd1 vccd1 vccd1 _16806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_234_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17786_ _17822_/CLK _17786_/D vssd1 vssd1 vccd1 vccd1 _17786_/Q sky130_fd_sc_hd__dfxtp_1
X_14998_ _15213_/A _15016_/B vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16737_ _17970_/CLK _16737_/D vssd1 vssd1 vccd1 vccd1 _16737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13949_ hold1271/X _13995_/A2 _13948_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _13949_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _18180_/CLK _16668_/D vssd1 vssd1 vccd1 vccd1 _16668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_232_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18407_ _18407_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_186_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15619_ _17269_/CLK _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _16631_/CLK _16599_/D vssd1 vssd1 vccd1 vccd1 _16599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09140_ _15523_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__or2_1
X_18338_ _18378_/CLK hold886/X vssd1 vssd1 vccd1 vccd1 hold885/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clkbuf_6_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09071_ hold1026/X _09119_/A2 _09070_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09071_/X
+ sky130_fd_sc_hd__o211a_1
X_18269_ _18409_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_272_wb_clk_i clkbuf_6_57_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08022_ hold1285/X _08029_/B _08021_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _08022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold701 hold701/A vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_201_wb_clk_i clkbuf_6_53_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18384_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold712 hold712/A vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold734 hold734/A vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold745 input59/X vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__clkbuf_2
Xhold756 hold756/A vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__buf_8
Xhold767 hold767/A vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold778 hold778/A vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ hold4777/X _10571_/B _09972_/X _15158_/C1 vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold789 hold789/A vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08924_ hold145/X hold156/X _08928_/S vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__mux2_1
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2102 _16169_/Q vssd1 vssd1 vccd1 vccd1 hold2102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2113 _17920_/Q vssd1 vssd1 vccd1 vccd1 hold2113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2124 hold2142/X vssd1 vssd1 vccd1 vccd1 hold2124/X sky130_fd_sc_hd__clkbuf_2
Xhold2135 _15550_/X vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 hold1401/A vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 _18298_/Q vssd1 vssd1 vccd1 vccd1 hold2146/X sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ _09053_/A hold307/X vssd1 vssd1 vccd1 vccd1 _16046_/D sky130_fd_sc_hd__and2_1
Xhold1412 _17750_/Q vssd1 vssd1 vccd1 vccd1 hold1412/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2157 _08008_/X vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2168 _15700_/Q vssd1 vssd1 vccd1 vccd1 hold2168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 _16183_/Q vssd1 vssd1 vccd1 vccd1 hold1423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 _16232_/Q vssd1 vssd1 vccd1 vccd1 hold2179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _15748_/Q vssd1 vssd1 vccd1 vccd1 hold1434/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1445 _07834_/X vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07806_ _07786_/A _07801_/B _09339_/B vssd1 vssd1 vccd1 vccd1 _07806_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1456 _15592_/Q vssd1 vssd1 vccd1 vccd1 hold1456/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1467 _15154_/X vssd1 vssd1 vccd1 vccd1 _18358_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ _15473_/A hold189/X vssd1 vssd1 vccd1 vccd1 _16013_/D sky130_fd_sc_hd__and2_1
Xhold1478 _08101_/X vssd1 vssd1 vccd1 vccd1 _15690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _15613_/Q vssd1 vssd1 vccd1 vccd1 hold1489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09407_ _07804_/A _09447_/C _15264_/A _09406_/X vssd1 vssd1 vccd1 vccd1 _09407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09338_ hold1897/X _09338_/A2 _09337_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _09338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09269_ hold181/X _16246_/Q _09273_/S vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11300_ _17770_/Q hold4662/X _12314_/C vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12280_ hold4273/X _12374_/B _12279_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ hold1173/X _16901_/Q _11711_/S vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ _16878_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__and3_1
XTAP_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4060 _09706_/X vssd1 vssd1 vccd1 vccd1 _16392_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _10497_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__or2_1
Xhold4071 _17182_/Q vssd1 vssd1 vccd1 vccd1 hold4071/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4082 _13336_/X vssd1 vssd1 vccd1 vccd1 _17565_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _18403_/CLK _15970_/D vssd1 vssd1 vccd1 vccd1 hold404/A sky130_fd_sc_hd__dfxtp_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ hold3088/X hold3914/X _11093_/S vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__mux2_1
Xhold4093 _17743_/Q vssd1 vssd1 vccd1 vccd1 hold4093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3370 _16485_/Q vssd1 vssd1 vccd1 vccd1 hold3370/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10044_ _13230_/A _09564_/A _10043_/X vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__a21oi_1
Xhold3381 _16421_/Q vssd1 vssd1 vccd1 vccd1 hold3381/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ hold3147/X _14952_/B _14920_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _14921_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3392 _16399_/Q vssd1 vssd1 vccd1 vccd1 hold3392/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__buf_6
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_6_18_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18040_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2680 _14925_/X vssd1 vssd1 vccd1 vccd1 _18247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _17738_/CLK _17640_/D vssd1 vssd1 vccd1 vccd1 _17640_/Q sky130_fd_sc_hd__dfxtp_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__buf_2
X_14852_ _15191_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__or2_1
XFILLER_0_216_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2691 _18394_/Q vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1990 _18175_/Q vssd1 vssd1 vccd1 vccd1 hold1990/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ hold3617/X _13713_/A _13802_/X vssd1 vssd1 vccd1 vccd1 _13803_/Y sky130_fd_sc_hd__a21oi_1
X_14783_ hold2353/X _14774_/B _14782_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14783_/X
+ sky130_fd_sc_hd__o211a_1
X_17571_ _17667_/CLK _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11995_ hold4382/X _13877_/B _11994_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_230_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16522_ _18078_/CLK _16522_/D vssd1 vssd1 vccd1 vccd1 _16522_/Q sky130_fd_sc_hd__dfxtp_1
X_13734_ _13734_/A _13734_/B vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10946_ hold1863/X _16806_/Q _11150_/C vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16453_ _18364_/CLK _16453_/D vssd1 vssd1 vccd1 vccd1 _16453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ _13761_/A _13665_/B vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__or2_1
X_10877_ hold645/X _16783_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15404_ _15482_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__and2_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ hold1261/X _17383_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16384_ _18327_/CLK _16384_/D vssd1 vssd1 vccd1 vccd1 _16384_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13788_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__or2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18123_ _18123_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
X_15335_ hold775/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12547_ hold2206/X hold3586/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15266_ _17330_/Q _15448_/B1 _09362_/D hold656/X vssd1 vssd1 vccd1 vccd1 _15266_/X
+ sky130_fd_sc_hd__a22o_1
X_18054_ _18054_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _17332_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14217_ _14897_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__or2_2
X_17005_ _17883_/CLK _17005_/D vssd1 vssd1 vccd1 vccd1 _17005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ hold3071/X _16967_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15197_ _15197_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _15547_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14079_ hold2409/X _14094_/B _14078_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__o211a_1
X_17907_ _17907_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_1
X_08640_ _12436_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _15942_/D sky130_fd_sc_hd__and2_1
X_17838_ _17891_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_238_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08571_ _12531_/A hold635/X vssd1 vssd1 vccd1 vccd1 _15909_/D sky130_fd_sc_hd__and2_1
X_17769_ _17769_/CLK _17769_/D vssd1 vssd1 vccd1 vccd1 hold697/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_453_wb_clk_i clkbuf_6_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09123_ _07788_/A _09120_/Y _09122_/Y _18457_/Q vssd1 vssd1 vccd1 vccd1 _09123_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ hold145/X hold424/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold425/A sky130_fd_sc_hd__mux2_1
XFILLER_0_142_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08005_ _14854_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold531 hold531/A vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__buf_2
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold553 input5/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold564 hold564/A vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold575 hold575/A vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 hold586/A vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold597/A vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09956_ hold1565/X hold3819/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08907_ _12424_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _16071_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ hold903/X hold3368/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__mux2_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _14559_/X vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 hold5827/X vssd1 vssd1 vccd1 vccd1 _13043_/C sky130_fd_sc_hd__buf_2
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ hold379/X hold827/X _08858_/S vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__mux2_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _08093_/X vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _09111_/X vssd1 vssd1 vccd1 vccd1 _16170_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 _14452_/X vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 la_data_in[12] vssd1 vssd1 vccd1 vccd1 hold1275/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1286 _08022_/X vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ hold402/X hold668/X _08779_/S vssd1 vssd1 vccd1 vccd1 hold669/A sky130_fd_sc_hd__mux2_1
Xhold1297 _09332_/X vssd1 vssd1 vccd1 vccd1 _16276_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _11121_/A _10800_/B vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__or2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11780_ _17084_/Q _12314_/B _12314_/C vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__and3_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _11667_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_194_wb_clk_i clkbuf_6_52_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ hold5739/X _13817_/B _13449_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10662_ _11052_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_123_wb_clk_i clkbuf_6_23_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12401_ hold98/X hold670/X _12401_/S vssd1 vssd1 vccd1 vccd1 hold671/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13381_ hold4583/X _13847_/B _13380_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10593_ hold3547/X _10497_/A _10592_/X vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15120_ hold2628/X _15111_/B _15119_/X _15198_/C1 vssd1 vssd1 vccd1 vccd1 _15120_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12332_ _17268_/Q _13868_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__and3_1
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15051_ _15105_/A hold2676/X _15071_/S vssd1 vssd1 vccd1 vccd1 _15052_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_239_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12263_ hold2212/X hold3470/X _13868_/C vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14002_ _14164_/A _14042_/B vssd1 vssd1 vccd1 vccd1 _14002_/X sky130_fd_sc_hd__or2_1
X_11214_ hold4693/X _11121_/A _11213_/X vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__a21oi_1
X_12194_ hold2302/X _17222_/Q _13412_/S vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput73 _13137_/A vssd1 vssd1 vccd1 vccd1 output73/X sky130_fd_sc_hd__buf_6
XFILLER_0_222_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ hold3679/X _11052_/A _11144_/X vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__a21oi_1
Xoutput84 _13217_/A vssd1 vssd1 vccd1 vccd1 output84/X sky130_fd_sc_hd__buf_6
XFILLER_0_222_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput95 _13297_/A vssd1 vssd1 vccd1 vccd1 output95/X sky130_fd_sc_hd__buf_6
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15953_ _17306_/CLK _15953_/D vssd1 vssd1 vccd1 vccd1 hold699/A sky130_fd_sc_hd__dfxtp_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11076_ _11643_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__or2_1
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ _11203_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _16499_/D sky130_fd_sc_hd__nor2_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14904_ _14974_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _17722_/CLK _15884_/D vssd1 vssd1 vccd1 vccd1 _15884_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _17623_/CLK _17623_/D vssd1 vssd1 vccd1 vccd1 _17623_/Q sky130_fd_sc_hd__dfxtp_1
X_14835_ hold3000/X _14826_/B _14834_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14835_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _18227_/CLK _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14766_ _15213_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__or2_1
X_11978_ hold1477/X _17150_/Q _12362_/C vssd1 vssd1 vccd1 vccd1 _11979_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16505_ _18384_/CLK _16505_/D vssd1 vssd1 vccd1 vccd1 _16505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _11121_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__or2_1
X_13717_ hold5030/X _13811_/B _13716_/X _08353_/A vssd1 vssd1 vccd1 vccd1 _13717_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_224_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14697_ hold1964/X _14720_/B _14696_/X _15222_/C1 vssd1 vssd1 vccd1 vccd1 _14697_/X
+ sky130_fd_sc_hd__o211a_1
X_17485_ _17485_/CLK _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16436_ _18379_/CLK _16436_/D vssd1 vssd1 vccd1 vccd1 _16436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ hold4309/X _13856_/B _13647_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13648_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _18342_/CLK _16367_/D vssd1 vssd1 vccd1 vccd1 _16367_/Q sky130_fd_sc_hd__dfxtp_1
X_13579_ hold5733/X _13817_/B _13578_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ _18170_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_1
X_15318_ hold405/X _15484_/A2 _09392_/D hold192/X vssd1 vssd1 vccd1 vccd1 _15318_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16298_ _16323_/CLK _16298_/D vssd1 vssd1 vccd1 vccd1 _16298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5508 _11500_/X vssd1 vssd1 vccd1 vccd1 _16990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5519 _16954_/Q vssd1 vssd1 vccd1 vccd1 hold5519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ _18071_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
X_15249_ hold326/X _15485_/A2 _15488_/A2 hold195/X _15248_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4807 _16884_/Q vssd1 vssd1 vccd1 vccd1 hold4807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4818 _09955_/X vssd1 vssd1 vccd1 vccd1 _16475_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4829 _16635_/Q vssd1 vssd1 vccd1 vccd1 hold4829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09810_ _09936_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__or2_1
Xfanout307 fanout334/X vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout318 _10527_/A vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__buf_4
Xfanout329 _09564_/A vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09741_ _09954_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__or2_1
XFILLER_0_201_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09672_ _09960_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_6_4_0_wb_clk_i clkbuf_6_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_6_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08623_ hold271/X hold308/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ hold361/X hold801/X _08592_/S vssd1 vssd1 vccd1 vccd1 hold802/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ hold2151/X _08488_/B _08484_/Y _08379_/A vssd1 vssd1 vccd1 vccd1 _08485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09106_ _15547_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_241_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09055_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _16135_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold361 hold23/X vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__clkbuf_8
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold394 hold394/A vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__buf_2
XFILLER_0_229_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout830 _14805_/C1 vssd1 vssd1 vccd1 vccd1 _14667_/C1 sky130_fd_sc_hd__buf_4
Xfanout841 _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14859_/C1 sky130_fd_sc_hd__buf_4
Xfanout852 _15217_/A vssd1 vssd1 vccd1 vccd1 _15543_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_217_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _09963_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__or2_1
Xfanout863 fanout873/X vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__buf_8
Xfanout874 hold819/X vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__buf_4
Xfanout885 _15195_/A vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__buf_8
X_12950_ hold3256/X _12949_/X _12998_/S vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__mux2_1
Xfanout896 _14116_/A vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__buf_8
XFILLER_0_232_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _16207_/Q vssd1 vssd1 vccd1 vccd1 hold1050/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1061 _15855_/Q vssd1 vssd1 vccd1 vccd1 hold1061/X sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _12024_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__or2_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1072 _18295_/Q vssd1 vssd1 vccd1 vccd1 hold1072/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 hold1134/X vssd1 vssd1 vccd1 vccd1 hold1135/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ hold3288/X _12880_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__mux2_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _18194_/Q vssd1 vssd1 vccd1 vccd1 hold1094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_375_wb_clk_i clkbuf_6_32_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17700_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14782_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14620_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11832_ _12261_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_304_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17896_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14551_ _15231_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__or2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ hold4815/X _11667_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ hold4887/X _11180_/B _10713_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__o211a_1
X_13502_ hold2053/X _17621_/Q _13874_/C vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__mux2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14482_ hold2701/X _14482_/A2 _14481_/Y _14542_/C1 vssd1 vssd1 vccd1 vccd1 _14482_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17270_/CLK _17270_/D vssd1 vssd1 vccd1 vccd1 _17270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11694_ _11694_/A _11694_/B vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13433_ _15835_/Q _17598_/Q _13817_/C vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__mux2_1
X_16221_ _17455_/CLK _16221_/D vssd1 vssd1 vccd1 vccd1 _16221_/Q sky130_fd_sc_hd__dfxtp_1
X_10645_ _11218_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _16705_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16152_ _17508_/CLK _16152_/D vssd1 vssd1 vccd1 vccd1 _16152_/Q sky130_fd_sc_hd__dfxtp_1
X_13364_ hold1687/X hold3328/X _13556_/S vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__mux2_1
X_10576_ _11194_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _16682_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15103_ _15103_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12315_ hold4653/X _12219_/A _12314_/X vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__a21oi_1
X_16083_ _16322_/CLK _16083_/D vssd1 vssd1 vccd1 vccd1 hold897/A sky130_fd_sc_hd__dfxtp_1
X_13295_ _13311_/A1 _13293_/X _13294_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15454_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__and2_1
X_12246_ _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_91_wb_clk_i clkbuf_6_17_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17286_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ _13782_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_6_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17459_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11128_ _11222_/A _11768_/B _11127_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11128_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16985_ _17863_/CLK _16985_/D vssd1 vssd1 vccd1 vccd1 _16985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15936_ _17326_/CLK _15936_/D vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__dfxtp_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _11153_/A _10019_/B _11058_/X _14434_/C1 vssd1 vssd1 vccd1 vccd1 _11059_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _17703_/CLK _15867_/D vssd1 vssd1 vccd1 vccd1 _15867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ _17702_/CLK _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14818_ _15211_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _17695_/CLK _15798_/D vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _18370_/CLK _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_1
X_14749_ hold2949/X _14772_/B _14748_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14749_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08270_ _15549_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17468_ _17469_/CLK _17468_/D vssd1 vssd1 vccd1 vccd1 _17468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16419_ _18266_/CLK _16419_/D vssd1 vssd1 vccd1 vccd1 _16419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ _18452_/CLK _17399_/D vssd1 vssd1 vccd1 vccd1 _17399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6006 data_in[24] vssd1 vssd1 vccd1 vccd1 hold575/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6017 la_data_in[21] vssd1 vssd1 vccd1 vccd1 hold556/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6028 data_in[10] vssd1 vssd1 vccd1 vccd1 hold570/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6039 _16523_/Q vssd1 vssd1 vccd1 vccd1 hold6039/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5305 _10891_/X vssd1 vssd1 vccd1 vccd1 _16787_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5316 _16589_/Q vssd1 vssd1 vccd1 vccd1 hold5316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5327 _11395_/X vssd1 vssd1 vccd1 vccd1 _16955_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5338 _17010_/Q vssd1 vssd1 vccd1 vccd1 hold5338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4604 _16352_/Q vssd1 vssd1 vccd1 vccd1 _13286_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5349 _11929_/X vssd1 vssd1 vccd1 vccd1 _17133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4615 _11181_/Y vssd1 vssd1 vccd1 vccd1 _11182_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4626 _11193_/Y vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4637 _16533_/Q vssd1 vssd1 vccd1 vccd1 hold4637/X sky130_fd_sc_hd__buf_1
XFILLER_0_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3903 _10150_/X vssd1 vssd1 vccd1 vccd1 _16540_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4648 _13812_/Y vssd1 vssd1 vccd1 vccd1 _13813_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3914 _16855_/Q vssd1 vssd1 vccd1 vccd1 hold3914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4659 _12306_/Y vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3925 _11248_/X vssd1 vssd1 vccd1 vccd1 _16906_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3936 _16469_/Q vssd1 vssd1 vccd1 vccd1 hold3936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3947 _09718_/X vssd1 vssd1 vccd1 vccd1 _16396_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3958 _16673_/Q vssd1 vssd1 vccd1 vccd1 hold3958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3969 _09508_/X vssd1 vssd1 vccd1 vccd1 _16326_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout148 _12755_/S vssd1 vssd1 vccd1 vccd1 _12773_/S sky130_fd_sc_hd__buf_6
Xfanout159 _12974_/S vssd1 vssd1 vccd1 vccd1 _12968_/S sky130_fd_sc_hd__buf_4
X_07985_ hold2717/X _07978_/B _07984_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09724_ hold5104/X _10010_/B _09723_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09724_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_236_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09655_ hold4763/X _10055_/B _09654_/X _15204_/C1 vssd1 vssd1 vccd1 vccd1 _09655_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08606_ _12426_/A _08606_/B vssd1 vssd1 vccd1 vccd1 _15925_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09586_ hold4731/X _10571_/B _09585_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09586_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ _09053_/A hold259/X vssd1 vssd1 vccd1 vccd1 _15892_/D sky130_fd_sc_hd__and2_1
XFILLER_0_132_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08468_ _14862_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08399_ _15513_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10430_ hold1829/X _16634_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ hold3086/X hold4805/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ hold5274/X _13798_/A2 _12099_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12100_/X
+ sky130_fd_sc_hd__o211a_1
X_13080_ _13073_/X _13079_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17528_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_131_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5850 hold5850/A vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_12
Xhold5861 _17522_/Q vssd1 vssd1 vccd1 vccd1 _13053_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_221_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10292_ hold1765/X _16588_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5872 hold5872/A vssd1 vssd1 vccd1 vccd1 hold5872/X sky130_fd_sc_hd__buf_2
Xhold5883 _16284_/Q vssd1 vssd1 vccd1 vccd1 hold5883/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12031_ hold4201/X _12031_/A2 _12030_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12031_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5894 hold5894/A vssd1 vssd1 vccd1 vccd1 hold5894/X sky130_fd_sc_hd__clkbuf_4
Xhold180 input46/X vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout660 _15502_/A vssd1 vssd1 vccd1 vccd1 _12894_/A sky130_fd_sc_hd__buf_4
Xfanout671 _08159_/A vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__buf_4
XFILLER_0_219_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout682 fanout692/X vssd1 vssd1 vccd1 vccd1 _15494_/A sky130_fd_sc_hd__clkbuf_4
X_16770_ _18003_/CLK _16770_/D vssd1 vssd1 vccd1 vccd1 _16770_/Q sky130_fd_sc_hd__dfxtp_1
X_13982_ _14878_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13982_/Y sky130_fd_sc_hd__nand2_1
Xfanout693 _07787_/Y vssd1 vssd1 vccd1 vccd1 fanout693/X sky130_fd_sc_hd__buf_4
XFILLER_0_219_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15721_ _17160_/CLK _15721_/D vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12999_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _17487_/D sky130_fd_sc_hd__and2_1
XFILLER_0_198_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18440_ _18442_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_35_0_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_6_35_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _17164_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12996_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _17464_/D sky130_fd_sc_hd__and2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ hold2405/X _14610_/B _14602_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14603_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18371_ _18371_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11815_ hold3812/X _12293_/B _11814_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _11815_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15583_ _17283_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12810_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _17441_/D sky130_fd_sc_hd__and2_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17322_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _17322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14534_ hold2909/X _14541_/B _14533_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14534_/X
+ sky130_fd_sc_hd__o211a_1
X_11746_ _13864_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _17072_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _17253_/CLK _17253_/D vssd1 vssd1 vccd1 vccd1 _17253_/Q sky130_fd_sc_hd__dfxtp_1
X_14465_ _14984_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__or2_1
X_11677_ hold5533/X _12338_/B _11676_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16204_ _17435_/CLK _16204_/D vssd1 vssd1 vccd1 vccd1 _16204_/Q sky130_fd_sc_hd__dfxtp_1
X_10628_ _16700_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10628_/X sky130_fd_sc_hd__and3_1
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13416_ _13800_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_226_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14396_ hold1837/X _14446_/A2 _14395_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17184_ _17280_/CLK _17184_/D vssd1 vssd1 vccd1 vccd1 _17184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16135_ _17330_/CLK _16135_/D vssd1 vssd1 vccd1 vccd1 hold632/A sky130_fd_sc_hd__dfxtp_1
X_13347_ _13767_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ hold1739/X _16677_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ _13278_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__or2_1
X_16066_ _17286_/CLK _16066_/D vssd1 vssd1 vccd1 vccd1 _16066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15017_ hold5982/X _15004_/B hold720/X _15162_/C1 vssd1 vssd1 vccd1 vccd1 hold721/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12229_ hold5489/X _12329_/B _12228_/X _08117_/A vssd1 vssd1 vccd1 vccd1 _12229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_227_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2509 _14143_/X vssd1 vssd1 vccd1 vccd1 _17873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1808 _15558_/X vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 _18360_/Q vssd1 vssd1 vccd1 vccd1 hold1819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_297_wb_clk_i clkbuf_6_39_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_237_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16968_ _17814_/CLK _16968_/D vssd1 vssd1 vccd1 vccd1 _16968_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_226_wb_clk_i clkbuf_6_61_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18213_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15919_ _18404_/CLK _15919_/D vssd1 vssd1 vccd1 vccd1 hold828/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16899_ _18068_/CLK _16899_/D vssd1 vssd1 vccd1 vccd1 _16899_/Q sky130_fd_sc_hd__dfxtp_1
X_09440_ _18462_/A _15304_/A vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__and2_1
XFILLER_0_232_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ hold433/X _15448_/B1 _15484_/B1 hold694/X _09370_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_75_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08322_ hold2451/X _08323_/B _08321_/Y _13720_/C1 vssd1 vssd1 vccd1 vccd1 _08322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08253_ hold2469/X _08263_/A2 _08252_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _08253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08184_ hold2100/X _08209_/B _08183_/X _08377_/A vssd1 vssd1 vccd1 vccd1 _08184_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5102 _16917_/Q vssd1 vssd1 vccd1 vccd1 hold5102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5113 _11092_/X vssd1 vssd1 vccd1 vccd1 _16854_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5124 _17020_/Q vssd1 vssd1 vccd1 vccd1 hold5124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5135 _11809_/X vssd1 vssd1 vccd1 vccd1 _17093_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5146 _17158_/Q vssd1 vssd1 vccd1 vccd1 hold5146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4401 _17185_/Q vssd1 vssd1 vccd1 vccd1 hold4401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4412 _12283_/X vssd1 vssd1 vccd1 vccd1 _17251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5157 _12013_/X vssd1 vssd1 vccd1 vccd1 _17161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5168 _16789_/Q vssd1 vssd1 vccd1 vccd1 hold5168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4423 _17247_/Q vssd1 vssd1 vccd1 vccd1 hold4423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4434 _11680_/X vssd1 vssd1 vccd1 vccd1 _17050_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5179 _10777_/X vssd1 vssd1 vccd1 vccd1 _16749_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3700 _13887_/Y vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4445 _17153_/Q vssd1 vssd1 vccd1 vccd1 hold4445/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3711 _10483_/X vssd1 vssd1 vccd1 vccd1 _16651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4456 _13567_/X vssd1 vssd1 vccd1 vccd1 _17642_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3722 _16922_/Q vssd1 vssd1 vccd1 vccd1 hold3722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4467 _16861_/Q vssd1 vssd1 vccd1 vccd1 hold4467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3733 _11142_/Y vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4478 _11983_/X vssd1 vssd1 vccd1 vccd1 _17151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3744 _16598_/Q vssd1 vssd1 vccd1 vccd1 hold3744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4489 _16873_/Q vssd1 vssd1 vccd1 vccd1 hold4489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3755 _10132_/X vssd1 vssd1 vccd1 vccd1 _16534_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3766 _16698_/Q vssd1 vssd1 vccd1 vccd1 hold3766/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3777 _10459_/X vssd1 vssd1 vccd1 vccd1 _16643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3788 _10432_/X vssd1 vssd1 vccd1 vccd1 _16634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3799 _17392_/Q vssd1 vssd1 vccd1 vccd1 hold3799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07968_ _15537_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09707_ hold2799/X _16393_/Q _10019_/C vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__mux2_1
X_07899_ hold2201/X _07918_/B _07898_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_223_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ hold1943/X hold5571/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ hold2490/X _16347_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ hold1610/X hold4293/X _12365_/C vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ hold2933/X _17371_/Q _12967_/S vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ hold2434/X hold3912/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14984_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11462_ hold2529/X hold5278/X _11738_/C vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _13201_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__and2_1
X_10413_ _10554_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10413_/X sky130_fd_sc_hd__or2_1
X_14181_ hold1973/X _14202_/B _14180_/X _13919_/A vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11393_ hold2804/X hold5320/X _12317_/C vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ hold4666/X _13131_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10344_ _10536_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5680 _09676_/X vssd1 vssd1 vccd1 vccd1 _16382_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13063_ _13199_/A1 _13061_/X _13062_/X _13199_/C1 vssd1 vssd1 vccd1 vccd1 _13063_/X
+ sky130_fd_sc_hd__o211a_2
X_17940_ _18035_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ _10563_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__or2_1
Xhold5691 _17709_/Q vssd1 vssd1 vccd1 vccd1 hold5691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12014_ hold2411/X hold4091/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__mux2_1
X_17871_ _17871_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4990 _16999_/Q vssd1 vssd1 vccd1 vccd1 hold4990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_390_wb_clk_i clkbuf_6_35_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16822_ _18055_/CLK _16822_/D vssd1 vssd1 vccd1 vccd1 _16822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout490 _10025_/C vssd1 vssd1 vccd1 vccd1 _11057_/S sky130_fd_sc_hd__buf_4
XFILLER_0_232_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16753_ _18018_/CLK _16753_/D vssd1 vssd1 vccd1 vccd1 _16753_/Q sky130_fd_sc_hd__dfxtp_1
X_13965_ hold3061/X _13995_/A2 _13964_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_232_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _17272_/CLK _15704_/D vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ hold2832/X _17483_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16684_ _18176_/CLK _16684_/D vssd1 vssd1 vccd1 vccd1 _16684_/Q sky130_fd_sc_hd__dfxtp_1
X_13896_ _15185_/A hold1501/X hold124/X vssd1 vssd1 vccd1 vccd1 _13896_/X sky130_fd_sc_hd__mux2_1
X_18423_ _18423_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15635_ _17179_/CLK _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ hold1464/X _17460_/Q _12913_/S vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18386_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _17234_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ hold2677/X hold3342/X _12808_/S vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17320_/CLK _17305_/D vssd1 vssd1 vccd1 vccd1 hold654/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _14517_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18285_ _18349_/CLK hold967/X vssd1 vssd1 vccd1 vccd1 hold966/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _17067_/Q _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__and3_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15497_ _14972_/A hold1544/X hold691/X vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _17236_/CLK _17236_/D vssd1 vssd1 vccd1 vccd1 _17236_/Q sky130_fd_sc_hd__dfxtp_1
X_14448_ _15128_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14479_/B sky130_fd_sc_hd__or2_4
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17167_ _17199_/CLK _17167_/D vssd1 vssd1 vccd1 vccd1 _17167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold905 hold905/A vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14379_ hold367/X hold658/X _14391_/S vssd1 vssd1 vccd1 vccd1 hold659/A sky130_fd_sc_hd__mux2_1
Xhold916 hold916/A vssd1 vssd1 vccd1 vccd1 hold916/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold927 hold927/A vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ _17346_/CLK _16118_/D vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__dfxtp_1
Xhold938 hold938/A vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 input68/X vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _17161_/CLK _17098_/D vssd1 vssd1 vccd1 vccd1 _17098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3007 _14707_/X vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16049_ _16097_/CLK _16049_/D vssd1 vssd1 vccd1 vccd1 hold304/A sky130_fd_sc_hd__dfxtp_1
X_08940_ _12412_/A hold884/X vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__and2_1
Xhold3018 _08247_/X vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3029 _18351_/Q vssd1 vssd1 vccd1 vccd1 hold3029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2306 _17811_/Q vssd1 vssd1 vccd1 vccd1 hold2306/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_407_wb_clk_i clkbuf_6_15_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17851_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08871_ _12386_/A hold662/X vssd1 vssd1 vccd1 vccd1 _16053_/D sky130_fd_sc_hd__and2_1
Xhold2317 _17922_/Q vssd1 vssd1 vccd1 vccd1 hold2317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2328 _08414_/X vssd1 vssd1 vccd1 vccd1 _15837_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2339 _18154_/Q vssd1 vssd1 vccd1 vccd1 hold2339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 _15763_/Q vssd1 vssd1 vccd1 vccd1 hold1605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ hold367/X hold181/A vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__or2_1
Xhold1616 _17896_/Q vssd1 vssd1 vccd1 vccd1 hold1616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1627 _14185_/X vssd1 vssd1 vccd1 vccd1 _17893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1638 _18270_/Q vssd1 vssd1 vccd1 vccd1 hold1638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 _15204_/X vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09423_ _07804_/A _09463_/A _15304_/A _09422_/X vssd1 vssd1 vccd1 vccd1 _09423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _09366_/A _09366_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09354_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_133_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08305_ _15203_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09285_ _14913_/A hold533/X vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08236_ _14116_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08167_ _08353_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08098_ _15557_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4220 _11044_/X vssd1 vssd1 vccd1 vccd1 _16838_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4231 _15998_/Q vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4242 _17407_/Q vssd1 vssd1 vccd1 vccd1 hold4242/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4253 _17188_/Q vssd1 vssd1 vccd1 vccd1 hold4253/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4264 _11965_/X vssd1 vssd1 vccd1 vccd1 _17145_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_148_wb_clk_i clkbuf_6_30_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18341_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3530 _13369_/X vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4275 _17004_/Q vssd1 vssd1 vccd1 vccd1 hold4275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _11194_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _16510_/D sky130_fd_sc_hd__nor2_1
Xhold3541 hold5843/X vssd1 vssd1 vccd1 vccd1 hold5844/A sky130_fd_sc_hd__buf_6
Xhold4286 _13471_/X vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3552 _10629_/Y vssd1 vssd1 vccd1 vccd1 _10630_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4297 _17648_/Q vssd1 vssd1 vccd1 vccd1 hold4297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3563 _16906_/Q vssd1 vssd1 vccd1 vccd1 hold3563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3574 _10005_/Y vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3585 _17368_/Q vssd1 vssd1 vccd1 vccd1 hold3585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2840 _18064_/Q vssd1 vssd1 vccd1 vccd1 hold2840/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2851 _14693_/X vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3596 _17113_/Q vssd1 vssd1 vccd1 vccd1 hold3596/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2862 _18188_/Q vssd1 vssd1 vccd1 vccd1 hold2862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2873 _07860_/X vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2884 _18091_/Q vssd1 vssd1 vccd1 vccd1 hold2884/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2895 _09099_/X vssd1 vssd1 vccd1 vccd1 _16164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10962_ _11136_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10962_/X sky130_fd_sc_hd__or2_1
X_13750_ hold3492/X _13883_/B _13749_/X _13750_/C1 vssd1 vssd1 vccd1 vccd1 _13750_/X
+ sky130_fd_sc_hd__o211a_1
X_12701_ hold3814/X _12700_/X _12764_/S vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _11082_/A _10893_/B vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__or2_1
X_13681_ hold4561/X _13777_/A2 _13680_/X _13777_/C1 vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15420_ hold298/X _09365_/B _09362_/D hold224/X _15418_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_183_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ hold3340/X _12631_/X _12809_/S vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ _16299_/Q _15477_/A2 _09392_/B hold883/X _15350_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/D sky130_fd_sc_hd__a221o_1
X_12563_ hold3599/X _12562_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14302_ _15523_/A _14336_/B vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__or2_1
X_11514_ _12246_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18070_ _18070_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
X_12494_ _17340_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__or2_1
X_15282_ _15489_/A _15282_/B _15282_/C _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_136_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17021_ _17804_/CLK _17021_/D vssd1 vssd1 vccd1 vccd1 _17021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11445_ _11637_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__or2_1
X_14233_ _14913_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14280_/B sky130_fd_sc_hd__or2_4
XFILLER_0_22_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14164_ _14164_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ _11694_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__or2_1
X_10327_ hold3950/X _10637_/B _10326_/X _14815_/C1 vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o211a_1
X_13115_ _13114_/X hold3600/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14095_ hold2510/X _14094_/B _14094_/Y _15496_/A vssd1 vssd1 vccd1 vccd1 _14095_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _17523_/Q hold960/X _13046_/C _13046_/D vssd1 vssd1 vccd1 vccd1 _13046_/X
+ sky130_fd_sc_hd__or4_1
X_17923_ _18018_/CLK _17923_/D vssd1 vssd1 vccd1 vccd1 _17923_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10258_ hold4164/X _10622_/B _10257_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17854_ _17886_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_1
X_10189_ hold5354/X _10625_/B _10188_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16805_ _18038_/CLK _16805_/D vssd1 vssd1 vccd1 vccd1 _16805_/Q sky130_fd_sc_hd__dfxtp_1
X_17785_ _18425_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
X_14997_ hold3015/X _15004_/B _14996_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _14997_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16736_ _18065_/CLK _16736_/D vssd1 vssd1 vccd1 vccd1 _16736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13948_ _15509_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16667_ _18223_/CLK _16667_/D vssd1 vssd1 vccd1 vccd1 _16667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ _13888_/A _13879_/B vssd1 vssd1 vccd1 vccd1 _17746_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_234_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18406_ _18406_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
X_15618_ _17234_/CLK _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16598_ _18198_/CLK _16598_/D vssd1 vssd1 vccd1 vccd1 _16598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ _18337_/CLK hold989/X vssd1 vssd1 vccd1 vccd1 hold988/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ _15549_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ hold999/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__or2_1
X_18268_ _18300_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _15535_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ _17283_/CLK _17219_/D vssd1 vssd1 vccd1 vccd1 _17219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18199_ _18199_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 hold724/A vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold735 hold735/A vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold746 hold746/A vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__buf_12
XFILLER_0_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold757 hold757/A vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 hold768/A vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _10470_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__or2_1
Xhold779 hold779/A vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_241_wb_clk_i clkbuf_6_62_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_228_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08923_ _15364_/A hold465/X vssd1 vssd1 vccd1 vccd1 _16079_/D sky130_fd_sc_hd__and2_1
Xhold2103 _09109_/X vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 _14243_/X vssd1 vssd1 vccd1 vccd1 _17920_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2125 _12512_/X vssd1 vssd1 vccd1 vccd1 _12974_/S sky130_fd_sc_hd__buf_4
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2136 _18437_/Q vssd1 vssd1 vccd1 vccd1 hold2136/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2147 _18050_/Q vssd1 vssd1 vccd1 vccd1 hold2147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 input38/X vssd1 vssd1 vccd1 vccd1 hold1402/X sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ hold222/X hold306/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1413 _07795_/X vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 _15839_/Q vssd1 vssd1 vccd1 vccd1 hold2158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 _09141_/X vssd1 vssd1 vccd1 vccd1 _16183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 _17759_/Q vssd1 vssd1 vccd1 vccd1 hold2169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_225_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1435 _08224_/X vssd1 vssd1 vccd1 vccd1 _15748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07805_/Y sky130_fd_sc_hd__inv_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1446 _17858_/Q vssd1 vssd1 vccd1 vccd1 hold1446/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08785_ hold145/X hold188/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__mux2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _07897_/X vssd1 vssd1 vccd1 vccd1 _15592_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _17890_/Q vssd1 vssd1 vccd1 vccd1 hold1468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_237_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1479 _18271_/Q vssd1 vssd1 vccd1 vccd1 hold1479/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09406_ _09438_/B _16289_/Q vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _15559_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _12747_/A hold105/X vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__and2_1
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08219_ _14726_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ hold991/X _09218_/B _09198_/X _12810_/A vssd1 vssd1 vccd1 vccd1 hold992/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_329_wb_clk_i clkbuf_6_44_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17904_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11230_ hold3829/X _11617_/A2 _11229_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11161_ _11203_/A _11161_/B vssd1 vssd1 vccd1 vccd1 _16877_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4050 _16492_/Q vssd1 vssd1 vccd1 vccd1 hold4050/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4061 _16659_/Q vssd1 vssd1 vccd1 vccd1 hold4061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ hold2703/X hold3547/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__mux2_1
XTAP_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4072 _11980_/X vssd1 vssd1 vccd1 vccd1 _17150_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ hold5112/X _11198_/B _11091_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _11092_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4083 _17656_/Q vssd1 vssd1 vccd1 vccd1 hold4083/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4094 _13774_/X vssd1 vssd1 vccd1 vccd1 _17711_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3360 _09643_/X vssd1 vssd1 vccd1 vccd1 _16371_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ _16505_/Q _10055_/B _10481_/S vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__and3_1
Xhold3371 _09889_/X vssd1 vssd1 vccd1 vccd1 _16453_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _15189_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__or2_1
Xhold3382 _09697_/X vssd1 vssd1 vccd1 vccd1 _16389_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3393 _09631_/X vssd1 vssd1 vccd1 vccd1 _16367_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__buf_6
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2670 _07862_/X vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ hold2989/X _14882_/B _14850_/X _14851_/C1 vssd1 vssd1 vccd1 vccd1 _14851_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2681 _18000_/Q vssd1 vssd1 vccd1 vccd1 hold2681/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_231_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2692 _15228_/X vssd1 vssd1 vccd1 vccd1 _18394_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13802_ _17721_/Q _13802_/B _13808_/C vssd1 vssd1 vccd1 vccd1 _13802_/X sky130_fd_sc_hd__and3_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _17730_/CLK _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1980 _08302_/X vssd1 vssd1 vccd1 vccd1 _15784_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1991 _14773_/X vssd1 vssd1 vccd1 vccd1 _18175_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _14782_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__or2_1
X_11994_ _13782_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__or2_1
X_16521_ _18233_/CLK _16521_/D vssd1 vssd1 vccd1 vccd1 _16521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ hold2557/X hold5701/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__mux2_1
X_10945_ hold5543/X _11156_/B _10944_/X _14366_/A vssd1 vssd1 vccd1 vccd1 _10945_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_230_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_wb_clk_i clkbuf_6_12_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _18395_/CLK _16452_/D vssd1 vssd1 vccd1 vccd1 _16452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13664_ hold2077/X _17675_/Q _13856_/C vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10876_ hold5559/X _11201_/B _10875_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _10876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15403_ _15481_/A1 _15395_/X _15402_/X _15481_/B1 hold5872/A vssd1 vssd1 vccd1 vccd1
+ _15403_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12615_ _12996_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _17381_/D sky130_fd_sc_hd__and2_1
X_16383_ _18294_/CLK _16383_/D vssd1 vssd1 vccd1 vccd1 _16383_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ hold2373/X hold4251/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13596_/B sky130_fd_sc_hd__mux2_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18122_ _18154_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15414_/A _15334_/B vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _12606_/A _12546_/B vssd1 vssd1 vccd1 vccd1 _17358_/D sky130_fd_sc_hd__and2_1
X_18053_ _18053_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
X_15265_ hold866/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15265_/X sky130_fd_sc_hd__or2_1
X_12477_ hold41/X _12445_/A _12445_/B _12476_/X _12436_/A vssd1 vssd1 vccd1 vccd1
+ hold42/A sky130_fd_sc_hd__o311a_1
XANTENNA_4 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _17882_/CLK _17004_/D vssd1 vssd1 vccd1 vccd1 _17004_/Q sky130_fd_sc_hd__dfxtp_1
X_14216_ _14897_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nor2_4
X_11428_ hold3772/X _12308_/B _11427_/X _15494_/A vssd1 vssd1 vccd1 vccd1 _11428_/X
+ sky130_fd_sc_hd__o211a_1
X_15196_ hold1054/X _15219_/B _15195_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14147_ hold2540/X _14148_/B _14146_/Y _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14147_/X
+ sky130_fd_sc_hd__o211a_1
X_11359_ hold4048/X _12314_/B _11358_/X _13927_/A vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14078_ _15531_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_238_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17906_ _17908_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_1
X_17837_ _17862_/CLK _17837_/D vssd1 vssd1 vccd1 vccd1 _17837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ hold402/X hold634/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold635/A sky130_fd_sc_hd__mux2_1
X_17768_ _17896_/CLK _17768_/D vssd1 vssd1 vccd1 vccd1 _17768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _17952_/CLK _16719_/D vssd1 vssd1 vccd1 vccd1 _16719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ _17731_/CLK _17699_/D vssd1 vssd1 vccd1 vccd1 _17699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09122_ _09122_/A _09122_/B vssd1 vssd1 vccd1 vccd1 _09122_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09053_ _09053_/A hold233/X vssd1 vssd1 vccd1 vccd1 _16143_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ hold2192/X _08033_/B _08003_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _08004_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_422_wb_clk_i clkbuf_6_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17200_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold510 hold749/X vssd1 vssd1 vccd1 vccd1 hold750/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_241_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold532 hold532/A vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold543 hold543/A vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold554 hold80/X vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__buf_4
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold58/X vssd1 vssd1 vccd1 vccd1 input21/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold587 hold587/A vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold598 hold598/A vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ hold4817/X _10049_/B _09954_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ hold568/X hold740/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__mux2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ hold5280/X _11159_/B _09885_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09886_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _17810_/Q vssd1 vssd1 vccd1 vccd1 hold1210/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _15614_/Q vssd1 vssd1 vccd1 vccd1 hold1221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 _18343_/Q vssd1 vssd1 vccd1 vccd1 hold1232/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _12416_/A _08837_/B vssd1 vssd1 vccd1 vccd1 _16037_/D sky130_fd_sc_hd__and2_1
Xhold1243 _15665_/Q vssd1 vssd1 vccd1 vccd1 hold1243/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1254 hold6036/X vssd1 vssd1 vccd1 vccd1 _09456_/C sky130_fd_sc_hd__clkbuf_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1265 _17800_/Q vssd1 vssd1 vccd1 vccd1 hold1265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 hold1276/A vssd1 vssd1 vccd1 vccd1 input40/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _17803_/Q vssd1 vssd1 vccd1 vccd1 hold1287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 _18215_/Q vssd1 vssd1 vccd1 vccd1 hold1298/X sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ _15394_/A hold569/X vssd1 vssd1 vccd1 vccd1 _16004_/D sky130_fd_sc_hd__and2_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08699_ hold379/X hold789/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10730_ hold2432/X hold4929/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10661_ hold1869/X hold3732/X _11147_/C vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _12408_/A hold321/X vssd1 vssd1 vccd1 vccd1 _17293_/D sky130_fd_sc_hd__and2_1
X_13380_ _13746_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10592_ _16688_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__and3_1
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12331_ _12340_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _17267_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_163_wb_clk_i clkbuf_6_27_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18397_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__and2_1
X_12262_ hold5421/X _13862_/B _12261_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12262_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11213_ _16895_/Q _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__and3_1
X_14001_ _14681_/A _14163_/B vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__or2_4
XFILLER_0_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ hold3821/X _13798_/A2 _12192_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11144_ _16872_/Q _11147_/B _11147_/C vssd1 vssd1 vccd1 vccd1 _11144_/X sky130_fd_sc_hd__and3_1
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput74 _13145_/A vssd1 vssd1 vccd1 vccd1 output74/X sky130_fd_sc_hd__buf_6
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 _13225_/A vssd1 vssd1 vccd1 vccd1 output85/X sky130_fd_sc_hd__buf_6
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 _13305_/A vssd1 vssd1 vccd1 vccd1 output96/X sky130_fd_sc_hd__buf_6
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _16087_/CLK _15952_/D vssd1 vssd1 vccd1 vccd1 hold909/A sky130_fd_sc_hd__dfxtp_1
X_11075_ hold2147/X _16849_/Q _11738_/C vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__mux2_1
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3190 _14593_/X vssd1 vssd1 vccd1 vccd1 _18088_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10026_ _13182_/A _11061_/A _10025_/X vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14903_ hold1805/X _14896_/Y _14902_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14903_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _17721_/CLK _15883_/D vssd1 vssd1 vccd1 vccd1 _15883_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _17686_/CLK _17622_/D vssd1 vssd1 vccd1 vccd1 _17622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14834_ _15227_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _18131_/CLK _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_230_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ hold3114/X _14772_/B _14764_/X _14835_/C1 vssd1 vssd1 vccd1 vccd1 _14765_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ hold3434/X _12347_/B _11976_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _18293_/CLK _16504_/D vssd1 vssd1 vccd1 vccd1 _16504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__or2_1
X_10928_ hold1697/X _16800_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__mux2_1
X_17484_ _17507_/CLK _17484_/D vssd1 vssd1 vccd1 vccd1 _17484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ _15197_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16435_ _18378_/CLK _16435_/D vssd1 vssd1 vccd1 vccd1 _16435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _13761_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__or2_1
X_10859_ hold2966/X _16777_/Q _11147_/C vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _18381_/CLK _16366_/D vssd1 vssd1 vccd1 vccd1 _16366_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13578_ _13698_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__or2_1
X_18105_ _18266_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ hold520/X _15487_/A2 _15484_/B1 hold415/X _15316_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12529_ hold1197/X _17354_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16297_ _17372_/CLK _16297_/D vssd1 vssd1 vccd1 vccd1 _16297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5509 _16946_/Q vssd1 vssd1 vccd1 vccd1 hold5509/X sky130_fd_sc_hd__dlygate4sd3_1
X_18036_ _18036_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ hold410/X _15484_/A2 _09392_/D hold340/X vssd1 vssd1 vccd1 vccd1 _15248_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4808 _11086_/X vssd1 vssd1 vccd1 vccd1 _16852_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4819 _16408_/Q vssd1 vssd1 vccd1 vccd1 hold4819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15179_ _15233_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout308 _11097_/A vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__buf_4
Xfanout319 _10527_/A vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__buf_4
XFILLER_0_158_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09740_ hold1178/X hold4743/X _10049_/C vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
.ends

