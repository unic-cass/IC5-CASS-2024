VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lovers_controller
  CLASS BLOCK ;
  FOREIGN lovers_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN becStatus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 546.000 74.890 550.000 ;
    END
  END becStatus[0]
  PIN becStatus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 546.000 81.790 550.000 ;
    END
  END becStatus[1]
  PIN becStatus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 546.000 88.690 550.000 ;
    END
  END becStatus[2]
  PIN becStatus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 95.310 546.000 95.590 550.000 ;
    END
  END becStatus[3]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 109.110 546.000 109.390 550.000 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 247.110 546.000 247.390 550.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 546.000 261.190 550.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 274.710 546.000 274.990 550.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 288.510 546.000 288.790 550.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 302.310 546.000 302.590 550.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 316.110 546.000 316.390 550.000 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 329.910 546.000 330.190 550.000 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 343.710 546.000 343.990 550.000 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 546.000 357.790 550.000 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 371.310 546.000 371.590 550.000 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 546.000 123.190 550.000 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 385.110 546.000 385.390 550.000 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 398.910 546.000 399.190 550.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 412.710 546.000 412.990 550.000 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 546.000 426.790 550.000 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 440.310 546.000 440.590 550.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 454.110 546.000 454.390 550.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 467.910 546.000 468.190 550.000 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 481.710 546.000 481.990 550.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 495.510 546.000 495.790 550.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 509.310 546.000 509.590 550.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 546.000 136.990 550.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 523.110 546.000 523.390 550.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 536.910 546.000 537.190 550.000 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 150.510 546.000 150.790 550.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 546.000 164.590 550.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 546.000 178.390 550.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 191.910 546.000 192.190 550.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 205.710 546.000 205.990 550.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.510 546.000 219.790 550.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 233.310 546.000 233.590 550.000 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 546.000 116.290 550.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 254.010 546.000 254.290 550.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 546.000 268.090 550.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 546.000 281.890 550.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 546.000 295.690 550.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 546.000 309.490 550.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 323.010 546.000 323.290 550.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 336.810 546.000 337.090 550.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 546.000 350.890 550.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 364.410 546.000 364.690 550.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 546.000 378.490 550.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 546.000 130.090 550.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.010 546.000 392.290 550.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 546.000 406.090 550.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 419.610 546.000 419.890 550.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 546.000 433.690 550.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 447.210 546.000 447.490 550.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 546.000 461.290 550.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 474.810 546.000 475.090 550.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 488.610 546.000 488.890 550.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 502.410 546.000 502.690 550.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 516.210 546.000 516.490 550.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 143.610 546.000 143.890 550.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 530.010 546.000 530.290 550.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 543.810 546.000 544.090 550.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 546.000 157.690 550.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 546.000 171.490 550.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 546.000 185.290 550.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 198.810 546.000 199.090 550.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 546.000 212.890 550.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 226.410 546.000 226.690 550.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 546.000 240.490 550.000 ;
    END
  END data_out[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 546.000 412.120 550.000 412.720 ;
    END
  END io_oeb
  PIN io_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 546.000 137.400 550.000 138.000 ;
    END
  END io_out
  PIN ki
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 546.000 54.190 550.000 ;
    END
  END ki
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END la_data_out[9]
  PIN load_data
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 546.000 47.290 550.000 ;
    END
  END load_data
  PIN load_status[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 5.610 546.000 5.890 550.000 ;
    END
  END load_status[0]
  PIN load_status[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 12.510 546.000 12.790 550.000 ;
    END
  END load_status[1]
  PIN load_status[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 546.000 19.690 550.000 ;
    END
  END load_status[2]
  PIN load_status[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 26.310 546.000 26.590 550.000 ;
    END
  END load_status[3]
  PIN load_status[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 546.000 33.490 550.000 ;
    END
  END load_status[4]
  PIN load_status[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 40.110 546.000 40.390 550.000 ;
    END
  END load_status[5]
  PIN next_key
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 60.810 546.000 61.090 550.000 ;
    END
  END next_key
  PIN slv_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 546.000 67.990 550.000 ;
    END
  END slv_done
  PIN slv_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 546.000 102.490 550.000 ;
    END
  END slv_enable
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 534.425 544.370 537.255 ;
        RECT 5.330 528.985 544.370 531.815 ;
        RECT 5.330 523.545 544.370 526.375 ;
        RECT 5.330 518.105 544.370 520.935 ;
        RECT 5.330 512.665 544.370 515.495 ;
        RECT 5.330 507.225 544.370 510.055 ;
        RECT 5.330 501.785 544.370 504.615 ;
        RECT 5.330 496.345 544.370 499.175 ;
        RECT 5.330 490.905 544.370 493.735 ;
        RECT 5.330 485.465 544.370 488.295 ;
        RECT 5.330 480.025 544.370 482.855 ;
        RECT 5.330 474.585 544.370 477.415 ;
        RECT 5.330 469.145 544.370 471.975 ;
        RECT 5.330 463.705 544.370 466.535 ;
        RECT 5.330 458.265 544.370 461.095 ;
        RECT 5.330 452.825 544.370 455.655 ;
        RECT 5.330 447.385 544.370 450.215 ;
        RECT 5.330 441.945 544.370 444.775 ;
        RECT 5.330 436.505 544.370 439.335 ;
        RECT 5.330 431.065 544.370 433.895 ;
        RECT 5.330 425.625 544.370 428.455 ;
        RECT 5.330 420.185 544.370 423.015 ;
        RECT 5.330 414.745 544.370 417.575 ;
        RECT 5.330 409.305 544.370 412.135 ;
        RECT 5.330 403.865 544.370 406.695 ;
        RECT 5.330 398.425 544.370 401.255 ;
        RECT 5.330 392.985 544.370 395.815 ;
        RECT 5.330 387.545 544.370 390.375 ;
        RECT 5.330 382.105 544.370 384.935 ;
        RECT 5.330 376.665 544.370 379.495 ;
        RECT 5.330 371.225 544.370 374.055 ;
        RECT 5.330 365.785 544.370 368.615 ;
        RECT 5.330 360.345 544.370 363.175 ;
        RECT 5.330 354.905 544.370 357.735 ;
        RECT 5.330 349.465 544.370 352.295 ;
        RECT 5.330 344.025 544.370 346.855 ;
        RECT 5.330 338.585 544.370 341.415 ;
        RECT 5.330 333.145 544.370 335.975 ;
        RECT 5.330 327.705 544.370 330.535 ;
        RECT 5.330 322.265 544.370 325.095 ;
        RECT 5.330 316.825 544.370 319.655 ;
        RECT 5.330 311.385 544.370 314.215 ;
        RECT 5.330 305.945 544.370 308.775 ;
        RECT 5.330 300.505 544.370 303.335 ;
        RECT 5.330 295.065 544.370 297.895 ;
        RECT 5.330 289.625 544.370 292.455 ;
        RECT 5.330 284.185 544.370 287.015 ;
        RECT 5.330 278.745 544.370 281.575 ;
        RECT 5.330 273.305 544.370 276.135 ;
        RECT 5.330 267.865 544.370 270.695 ;
        RECT 5.330 262.425 544.370 265.255 ;
        RECT 5.330 256.985 544.370 259.815 ;
        RECT 5.330 251.545 544.370 254.375 ;
        RECT 5.330 246.105 544.370 248.935 ;
        RECT 5.330 240.665 544.370 243.495 ;
        RECT 5.330 235.225 544.370 238.055 ;
        RECT 5.330 229.785 544.370 232.615 ;
        RECT 5.330 224.345 544.370 227.175 ;
        RECT 5.330 218.905 544.370 221.735 ;
        RECT 5.330 213.465 544.370 216.295 ;
        RECT 5.330 208.025 544.370 210.855 ;
        RECT 5.330 202.585 544.370 205.415 ;
        RECT 5.330 197.145 544.370 199.975 ;
        RECT 5.330 191.705 544.370 194.535 ;
        RECT 5.330 186.265 544.370 189.095 ;
        RECT 5.330 180.825 544.370 183.655 ;
        RECT 5.330 175.385 544.370 178.215 ;
        RECT 5.330 169.945 544.370 172.775 ;
        RECT 5.330 164.505 544.370 167.335 ;
        RECT 5.330 159.065 544.370 161.895 ;
        RECT 5.330 153.625 544.370 156.455 ;
        RECT 5.330 148.185 544.370 151.015 ;
        RECT 5.330 142.745 544.370 145.575 ;
        RECT 5.330 137.305 544.370 140.135 ;
        RECT 5.330 131.865 544.370 134.695 ;
        RECT 5.330 126.425 544.370 129.255 ;
        RECT 5.330 120.985 544.370 123.815 ;
        RECT 5.330 115.545 544.370 118.375 ;
        RECT 5.330 110.105 544.370 112.935 ;
        RECT 5.330 104.665 544.370 107.495 ;
        RECT 5.330 99.225 544.370 102.055 ;
        RECT 5.330 93.785 544.370 96.615 ;
        RECT 5.330 88.345 544.370 91.175 ;
        RECT 5.330 82.905 544.370 85.735 ;
        RECT 5.330 77.465 544.370 80.295 ;
        RECT 5.330 72.025 544.370 74.855 ;
        RECT 5.330 66.585 544.370 69.415 ;
        RECT 5.330 61.145 544.370 63.975 ;
        RECT 5.330 55.705 544.370 58.535 ;
        RECT 5.330 50.265 544.370 53.095 ;
        RECT 5.330 44.825 544.370 47.655 ;
        RECT 5.330 39.385 544.370 42.215 ;
        RECT 5.330 33.945 544.370 36.775 ;
        RECT 5.330 28.505 544.370 31.335 ;
        RECT 5.330 23.065 544.370 25.895 ;
        RECT 5.330 17.625 544.370 20.455 ;
        RECT 5.330 12.185 544.370 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 5.520 7.180 544.480 540.560 ;
      LAYER met2 ;
        RECT 6.170 545.720 12.230 546.450 ;
        RECT 13.070 545.720 19.130 546.450 ;
        RECT 19.970 545.720 26.030 546.450 ;
        RECT 26.870 545.720 32.930 546.450 ;
        RECT 33.770 545.720 39.830 546.450 ;
        RECT 40.670 545.720 46.730 546.450 ;
        RECT 47.570 545.720 53.630 546.450 ;
        RECT 54.470 545.720 60.530 546.450 ;
        RECT 61.370 545.720 67.430 546.450 ;
        RECT 68.270 545.720 74.330 546.450 ;
        RECT 75.170 545.720 81.230 546.450 ;
        RECT 82.070 545.720 88.130 546.450 ;
        RECT 88.970 545.720 95.030 546.450 ;
        RECT 95.870 545.720 101.930 546.450 ;
        RECT 102.770 545.720 108.830 546.450 ;
        RECT 109.670 545.720 115.730 546.450 ;
        RECT 116.570 545.720 122.630 546.450 ;
        RECT 123.470 545.720 129.530 546.450 ;
        RECT 130.370 545.720 136.430 546.450 ;
        RECT 137.270 545.720 143.330 546.450 ;
        RECT 144.170 545.720 150.230 546.450 ;
        RECT 151.070 545.720 157.130 546.450 ;
        RECT 157.970 545.720 164.030 546.450 ;
        RECT 164.870 545.720 170.930 546.450 ;
        RECT 171.770 545.720 177.830 546.450 ;
        RECT 178.670 545.720 184.730 546.450 ;
        RECT 185.570 545.720 191.630 546.450 ;
        RECT 192.470 545.720 198.530 546.450 ;
        RECT 199.370 545.720 205.430 546.450 ;
        RECT 206.270 545.720 212.330 546.450 ;
        RECT 213.170 545.720 219.230 546.450 ;
        RECT 220.070 545.720 226.130 546.450 ;
        RECT 226.970 545.720 233.030 546.450 ;
        RECT 233.870 545.720 239.930 546.450 ;
        RECT 240.770 545.720 246.830 546.450 ;
        RECT 247.670 545.720 253.730 546.450 ;
        RECT 254.570 545.720 260.630 546.450 ;
        RECT 261.470 545.720 267.530 546.450 ;
        RECT 268.370 545.720 274.430 546.450 ;
        RECT 275.270 545.720 281.330 546.450 ;
        RECT 282.170 545.720 288.230 546.450 ;
        RECT 289.070 545.720 295.130 546.450 ;
        RECT 295.970 545.720 302.030 546.450 ;
        RECT 302.870 545.720 308.930 546.450 ;
        RECT 309.770 545.720 315.830 546.450 ;
        RECT 316.670 545.720 322.730 546.450 ;
        RECT 323.570 545.720 329.630 546.450 ;
        RECT 330.470 545.720 336.530 546.450 ;
        RECT 337.370 545.720 343.430 546.450 ;
        RECT 344.270 545.720 350.330 546.450 ;
        RECT 351.170 545.720 357.230 546.450 ;
        RECT 358.070 545.720 364.130 546.450 ;
        RECT 364.970 545.720 371.030 546.450 ;
        RECT 371.870 545.720 377.930 546.450 ;
        RECT 378.770 545.720 384.830 546.450 ;
        RECT 385.670 545.720 391.730 546.450 ;
        RECT 392.570 545.720 398.630 546.450 ;
        RECT 399.470 545.720 405.530 546.450 ;
        RECT 406.370 545.720 412.430 546.450 ;
        RECT 413.270 545.720 419.330 546.450 ;
        RECT 420.170 545.720 426.230 546.450 ;
        RECT 427.070 545.720 433.130 546.450 ;
        RECT 433.970 545.720 440.030 546.450 ;
        RECT 440.870 545.720 446.930 546.450 ;
        RECT 447.770 545.720 453.830 546.450 ;
        RECT 454.670 545.720 460.730 546.450 ;
        RECT 461.570 545.720 467.630 546.450 ;
        RECT 468.470 545.720 474.530 546.450 ;
        RECT 475.370 545.720 481.430 546.450 ;
        RECT 482.270 545.720 488.330 546.450 ;
        RECT 489.170 545.720 495.230 546.450 ;
        RECT 496.070 545.720 502.130 546.450 ;
        RECT 502.970 545.720 509.030 546.450 ;
        RECT 509.870 545.720 515.930 546.450 ;
        RECT 516.770 545.720 522.830 546.450 ;
        RECT 523.670 545.720 529.730 546.450 ;
        RECT 530.570 545.720 536.630 546.450 ;
        RECT 537.470 545.720 543.530 546.450 ;
        RECT 5.620 4.280 544.080 545.720 ;
        RECT 6.170 3.670 13.610 4.280 ;
        RECT 14.450 3.670 21.890 4.280 ;
        RECT 22.730 3.670 30.170 4.280 ;
        RECT 31.010 3.670 38.450 4.280 ;
        RECT 39.290 3.670 46.730 4.280 ;
        RECT 47.570 3.670 55.010 4.280 ;
        RECT 55.850 3.670 63.290 4.280 ;
        RECT 64.130 3.670 71.570 4.280 ;
        RECT 72.410 3.670 79.850 4.280 ;
        RECT 80.690 3.670 88.130 4.280 ;
        RECT 88.970 3.670 96.410 4.280 ;
        RECT 97.250 3.670 104.690 4.280 ;
        RECT 105.530 3.670 112.970 4.280 ;
        RECT 113.810 3.670 121.250 4.280 ;
        RECT 122.090 3.670 129.530 4.280 ;
        RECT 130.370 3.670 137.810 4.280 ;
        RECT 138.650 3.670 146.090 4.280 ;
        RECT 146.930 3.670 154.370 4.280 ;
        RECT 155.210 3.670 162.650 4.280 ;
        RECT 163.490 3.670 170.930 4.280 ;
        RECT 171.770 3.670 179.210 4.280 ;
        RECT 180.050 3.670 187.490 4.280 ;
        RECT 188.330 3.670 195.770 4.280 ;
        RECT 196.610 3.670 204.050 4.280 ;
        RECT 204.890 3.670 212.330 4.280 ;
        RECT 213.170 3.670 220.610 4.280 ;
        RECT 221.450 3.670 228.890 4.280 ;
        RECT 229.730 3.670 237.170 4.280 ;
        RECT 238.010 3.670 245.450 4.280 ;
        RECT 246.290 3.670 253.730 4.280 ;
        RECT 254.570 3.670 262.010 4.280 ;
        RECT 262.850 3.670 270.290 4.280 ;
        RECT 271.130 3.670 278.570 4.280 ;
        RECT 279.410 3.670 286.850 4.280 ;
        RECT 287.690 3.670 295.130 4.280 ;
        RECT 295.970 3.670 303.410 4.280 ;
        RECT 304.250 3.670 311.690 4.280 ;
        RECT 312.530 3.670 319.970 4.280 ;
        RECT 320.810 3.670 328.250 4.280 ;
        RECT 329.090 3.670 336.530 4.280 ;
        RECT 337.370 3.670 344.810 4.280 ;
        RECT 345.650 3.670 353.090 4.280 ;
        RECT 353.930 3.670 361.370 4.280 ;
        RECT 362.210 3.670 369.650 4.280 ;
        RECT 370.490 3.670 377.930 4.280 ;
        RECT 378.770 3.670 386.210 4.280 ;
        RECT 387.050 3.670 394.490 4.280 ;
        RECT 395.330 3.670 402.770 4.280 ;
        RECT 403.610 3.670 411.050 4.280 ;
        RECT 411.890 3.670 419.330 4.280 ;
        RECT 420.170 3.670 427.610 4.280 ;
        RECT 428.450 3.670 435.890 4.280 ;
        RECT 436.730 3.670 444.170 4.280 ;
        RECT 445.010 3.670 452.450 4.280 ;
        RECT 453.290 3.670 460.730 4.280 ;
        RECT 461.570 3.670 469.010 4.280 ;
        RECT 469.850 3.670 477.290 4.280 ;
        RECT 478.130 3.670 485.570 4.280 ;
        RECT 486.410 3.670 493.850 4.280 ;
        RECT 494.690 3.670 502.130 4.280 ;
        RECT 502.970 3.670 510.410 4.280 ;
        RECT 511.250 3.670 518.690 4.280 ;
        RECT 519.530 3.670 526.970 4.280 ;
        RECT 527.810 3.670 535.250 4.280 ;
        RECT 536.090 3.670 543.530 4.280 ;
      LAYER met3 ;
        RECT 20.305 413.120 546.000 540.425 ;
        RECT 20.305 411.720 545.600 413.120 ;
        RECT 20.305 138.400 546.000 411.720 ;
        RECT 20.305 137.000 545.600 138.400 ;
        RECT 20.305 8.335 546.000 137.000 ;
      LAYER met4 ;
        RECT 23.295 539.200 513.065 540.425 ;
        RECT 23.295 10.240 97.440 539.200 ;
        RECT 99.840 10.240 174.240 539.200 ;
        RECT 176.640 10.240 251.040 539.200 ;
        RECT 253.440 10.240 327.840 539.200 ;
        RECT 330.240 10.240 404.640 539.200 ;
        RECT 407.040 10.240 481.440 539.200 ;
        RECT 483.840 10.240 513.065 539.200 ;
        RECT 23.295 8.335 513.065 10.240 ;
  END
END lovers_controller
END LIBRARY

