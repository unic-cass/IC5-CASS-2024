magic
tech sky130A
magscale 1 2
timestamp 1731520197
<< obsli1 >>
rect 1104 2159 158884 127313
<< obsm1 >>
rect 198 76 159882 127344
<< metal2 >>
rect 2686 0 2742 800
rect 4618 0 4674 800
rect 6550 0 6606 800
rect 8482 0 8538 800
rect 10414 0 10470 800
rect 12346 0 12402 800
rect 14278 0 14334 800
rect 16210 0 16266 800
rect 18142 0 18198 800
rect 20074 0 20130 800
rect 22006 0 22062 800
rect 23938 0 23994 800
rect 25870 0 25926 800
rect 27802 0 27858 800
rect 29734 0 29790 800
rect 31666 0 31722 800
rect 33598 0 33654 800
rect 35530 0 35586 800
rect 37462 0 37518 800
rect 39394 0 39450 800
rect 41326 0 41382 800
rect 43258 0 43314 800
rect 45190 0 45246 800
rect 47122 0 47178 800
rect 49054 0 49110 800
rect 50986 0 51042 800
rect 52918 0 52974 800
rect 54850 0 54906 800
rect 56782 0 56838 800
rect 58714 0 58770 800
rect 60646 0 60702 800
rect 62578 0 62634 800
rect 64510 0 64566 800
rect 66442 0 66498 800
rect 68374 0 68430 800
rect 70306 0 70362 800
rect 72238 0 72294 800
rect 74170 0 74226 800
rect 76102 0 76158 800
rect 78034 0 78090 800
rect 79966 0 80022 800
rect 81898 0 81954 800
rect 83830 0 83886 800
rect 85762 0 85818 800
rect 87694 0 87750 800
rect 89626 0 89682 800
rect 91558 0 91614 800
rect 93490 0 93546 800
rect 95422 0 95478 800
rect 97354 0 97410 800
rect 99286 0 99342 800
rect 101218 0 101274 800
rect 103150 0 103206 800
rect 105082 0 105138 800
rect 107014 0 107070 800
rect 108946 0 109002 800
rect 110878 0 110934 800
rect 112810 0 112866 800
rect 114742 0 114798 800
rect 116674 0 116730 800
rect 118606 0 118662 800
rect 120538 0 120594 800
rect 122470 0 122526 800
rect 124402 0 124458 800
rect 126334 0 126390 800
rect 128266 0 128322 800
rect 130198 0 130254 800
rect 132130 0 132186 800
rect 134062 0 134118 800
rect 135994 0 136050 800
rect 137926 0 137982 800
rect 139858 0 139914 800
rect 141790 0 141846 800
rect 143722 0 143778 800
rect 145654 0 145710 800
rect 147586 0 147642 800
rect 149518 0 149574 800
rect 151450 0 151506 800
rect 153382 0 153438 800
rect 155314 0 155370 800
rect 157246 0 157302 800
<< obsm2 >>
rect 204 856 159876 127333
rect 204 31 2630 856
rect 2798 31 4562 856
rect 4730 31 6494 856
rect 6662 31 8426 856
rect 8594 31 10358 856
rect 10526 31 12290 856
rect 12458 31 14222 856
rect 14390 31 16154 856
rect 16322 31 18086 856
rect 18254 31 20018 856
rect 20186 31 21950 856
rect 22118 31 23882 856
rect 24050 31 25814 856
rect 25982 31 27746 856
rect 27914 31 29678 856
rect 29846 31 31610 856
rect 31778 31 33542 856
rect 33710 31 35474 856
rect 35642 31 37406 856
rect 37574 31 39338 856
rect 39506 31 41270 856
rect 41438 31 43202 856
rect 43370 31 45134 856
rect 45302 31 47066 856
rect 47234 31 48998 856
rect 49166 31 50930 856
rect 51098 31 52862 856
rect 53030 31 54794 856
rect 54962 31 56726 856
rect 56894 31 58658 856
rect 58826 31 60590 856
rect 60758 31 62522 856
rect 62690 31 64454 856
rect 64622 31 66386 856
rect 66554 31 68318 856
rect 68486 31 70250 856
rect 70418 31 72182 856
rect 72350 31 74114 856
rect 74282 31 76046 856
rect 76214 31 77978 856
rect 78146 31 79910 856
rect 80078 31 81842 856
rect 82010 31 83774 856
rect 83942 31 85706 856
rect 85874 31 87638 856
rect 87806 31 89570 856
rect 89738 31 91502 856
rect 91670 31 93434 856
rect 93602 31 95366 856
rect 95534 31 97298 856
rect 97466 31 99230 856
rect 99398 31 101162 856
rect 101330 31 103094 856
rect 103262 31 105026 856
rect 105194 31 106958 856
rect 107126 31 108890 856
rect 109058 31 110822 856
rect 110990 31 112754 856
rect 112922 31 114686 856
rect 114854 31 116618 856
rect 116786 31 118550 856
rect 118718 31 120482 856
rect 120650 31 122414 856
rect 122582 31 124346 856
rect 124514 31 126278 856
rect 126446 31 128210 856
rect 128378 31 130142 856
rect 130310 31 132074 856
rect 132242 31 134006 856
rect 134174 31 135938 856
rect 136106 31 137870 856
rect 138038 31 139802 856
rect 139970 31 141734 856
rect 141902 31 143666 856
rect 143834 31 145598 856
rect 145766 31 147530 856
rect 147698 31 149462 856
rect 149630 31 151394 856
rect 151562 31 153326 856
rect 153494 31 155258 856
rect 155426 31 157190 856
rect 157358 31 159876 856
<< obsm3 >>
rect 289 35 159791 127329
<< metal4 >>
rect 4208 2128 4528 127344
rect 19568 2128 19888 127344
rect 34928 2128 35248 127344
rect 50288 2128 50608 127344
rect 65648 2128 65968 127344
rect 81008 2128 81328 127344
rect 96368 2128 96688 127344
rect 111728 2128 112048 127344
rect 127088 2128 127408 127344
rect 142448 2128 142768 127344
rect 157808 2128 158128 127344
<< obsm4 >>
rect 427 2048 4128 121549
rect 4608 2048 19488 121549
rect 19968 2048 34848 121549
rect 35328 2048 50208 121549
rect 50688 2048 65568 121549
rect 66048 2048 80928 121549
rect 81408 2048 96288 121549
rect 96768 2048 111648 121549
rect 112128 2048 127008 121549
rect 127488 2048 142368 121549
rect 142848 2048 157445 121549
rect 427 443 157445 2048
<< labels >>
rlabel metal2 s 27802 0 27858 800 6 becStatus[0]
port 1 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 becStatus[1]
port 2 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 becStatus[2]
port 3 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 becStatus[3]
port 4 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 clk
port 5 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 data_in[0]
port 6 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 data_in[10]
port 7 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 data_in[11]
port 8 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 data_in[12]
port 9 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 data_in[13]
port 10 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 data_in[14]
port 11 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 data_in[15]
port 12 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 data_in[16]
port 13 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 data_in[17]
port 14 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 data_in[18]
port 15 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 data_in[19]
port 16 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 data_in[1]
port 17 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 data_in[20]
port 18 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 data_in[21]
port 19 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 data_in[22]
port 20 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 data_in[23]
port 21 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 data_in[24]
port 22 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 data_in[25]
port 23 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 data_in[26]
port 24 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 data_in[27]
port 25 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 data_in[28]
port 26 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 data_in[29]
port 27 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 data_in[2]
port 28 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 data_in[30]
port 29 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 data_in[31]
port 30 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 data_in[3]
port 31 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 data_in[4]
port 32 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 data_in[5]
port 33 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 data_in[6]
port 34 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 data_in[7]
port 35 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 data_in[8]
port 36 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 data_in[9]
port 37 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 data_out[0]
port 38 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 data_out[10]
port 39 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 data_out[11]
port 40 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 data_out[12]
port 41 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 data_out[13]
port 42 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 data_out[14]
port 43 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 data_out[15]
port 44 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 data_out[16]
port 45 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 data_out[17]
port 46 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 data_out[18]
port 47 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 data_out[19]
port 48 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 data_out[1]
port 49 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 data_out[20]
port 50 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 data_out[21]
port 51 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 data_out[22]
port 52 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 data_out[23]
port 53 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 data_out[24]
port 54 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 data_out[25]
port 55 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 data_out[26]
port 56 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 data_out[27]
port 57 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 data_out[28]
port 58 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 data_out[29]
port 59 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 data_out[2]
port 60 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 data_out[30]
port 61 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 data_out[31]
port 62 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 data_out[3]
port 63 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 data_out[4]
port 64 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 data_out[5]
port 65 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 data_out[6]
port 66 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 data_out[7]
port 67 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 data_out[8]
port 68 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 data_out[9]
port 69 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 done
port 70 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 enable
port 71 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 ki
port 72 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 load_data
port 73 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 load_status[0]
port 74 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 load_status[1]
port 75 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 load_status[2]
port 76 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 load_status[3]
port 77 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 load_status[4]
port 78 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 load_status[5]
port 79 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 next_key
port 80 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 rst
port 81 nsew signal input
rlabel metal4 s 4208 2128 4528 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 127344 6 vccd2
port 82 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 127344 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 127344 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 127344 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 127344 6 vssd2
port 83 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 127344 6 vssd2
port 83 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 160000 130000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 64672088
string GDS_FILE /home/cass/projects/IC5-CASS-2024/openlane/lovers_bec/runs/24_11_13_23_48/results/signoff/bec.magic.gds
string GDS_START 881448
<< end >>

