VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc_wrapper
  CLASS BLOCK ;
  FOREIGN vco_adc_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1264.440 BY 1275.160 ;
  PIN phase_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 316.110 1271.160 316.390 1275.160 ;
    END
  END phase_in
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1262.320 ;
    END
  END vccd1
  PIN vco_enb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 948.150 1271.160 948.430 1275.160 ;
    END
  END vco_enb_o
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1262.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1262.320 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1005.650 0.000 1005.930 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 0.000 1189.930 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 925.150 0.000 925.430 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1132.150 0.000 1132.430 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 1257.945 1258.750 1260.775 ;
        RECT 5.330 1252.505 1258.750 1255.335 ;
        RECT 5.330 1247.065 1258.750 1249.895 ;
        RECT 5.330 1241.625 1258.750 1244.455 ;
        RECT 5.330 1236.185 1258.750 1239.015 ;
        RECT 5.330 1230.745 1258.750 1233.575 ;
        RECT 5.330 1225.305 1258.750 1228.135 ;
        RECT 5.330 1219.865 1258.750 1222.695 ;
        RECT 5.330 1214.425 1258.750 1217.255 ;
        RECT 5.330 1208.985 1258.750 1211.815 ;
        RECT 5.330 1203.545 1258.750 1206.375 ;
        RECT 5.330 1198.105 1258.750 1200.935 ;
        RECT 5.330 1192.665 1258.750 1195.495 ;
        RECT 5.330 1187.225 1258.750 1190.055 ;
        RECT 5.330 1181.785 1258.750 1184.615 ;
        RECT 5.330 1176.345 1258.750 1179.175 ;
        RECT 5.330 1170.905 1258.750 1173.735 ;
        RECT 5.330 1165.465 1258.750 1168.295 ;
        RECT 5.330 1160.025 1258.750 1162.855 ;
        RECT 5.330 1154.585 1258.750 1157.415 ;
        RECT 5.330 1149.145 1258.750 1151.975 ;
        RECT 5.330 1143.705 1258.750 1146.535 ;
        RECT 5.330 1138.265 1258.750 1141.095 ;
        RECT 5.330 1132.825 1258.750 1135.655 ;
        RECT 5.330 1127.385 1258.750 1130.215 ;
        RECT 5.330 1121.945 1258.750 1124.775 ;
        RECT 5.330 1116.505 1258.750 1119.335 ;
        RECT 5.330 1111.065 1258.750 1113.895 ;
        RECT 5.330 1105.625 1258.750 1108.455 ;
        RECT 5.330 1100.185 1258.750 1103.015 ;
        RECT 5.330 1094.745 1258.750 1097.575 ;
        RECT 5.330 1089.305 1258.750 1092.135 ;
        RECT 5.330 1083.865 1258.750 1086.695 ;
        RECT 5.330 1078.425 1258.750 1081.255 ;
        RECT 5.330 1072.985 1258.750 1075.815 ;
        RECT 5.330 1067.545 1258.750 1070.375 ;
        RECT 5.330 1062.105 1258.750 1064.935 ;
        RECT 5.330 1056.665 1258.750 1059.495 ;
        RECT 5.330 1051.225 1258.750 1054.055 ;
        RECT 5.330 1045.785 1258.750 1048.615 ;
        RECT 5.330 1040.345 1258.750 1043.175 ;
        RECT 5.330 1034.905 1258.750 1037.735 ;
        RECT 5.330 1029.465 1258.750 1032.295 ;
        RECT 5.330 1024.025 1258.750 1026.855 ;
        RECT 5.330 1018.585 1258.750 1021.415 ;
        RECT 5.330 1013.145 1258.750 1015.975 ;
        RECT 5.330 1007.705 1258.750 1010.535 ;
        RECT 5.330 1002.265 1258.750 1005.095 ;
        RECT 5.330 996.825 1258.750 999.655 ;
        RECT 5.330 991.385 1258.750 994.215 ;
        RECT 5.330 985.945 1258.750 988.775 ;
        RECT 5.330 980.505 1258.750 983.335 ;
        RECT 5.330 975.065 1258.750 977.895 ;
        RECT 5.330 969.625 1258.750 972.455 ;
        RECT 5.330 964.185 1258.750 967.015 ;
        RECT 5.330 958.745 1258.750 961.575 ;
        RECT 5.330 953.305 1258.750 956.135 ;
        RECT 5.330 947.865 1258.750 950.695 ;
        RECT 5.330 942.425 1258.750 945.255 ;
        RECT 5.330 936.985 1258.750 939.815 ;
        RECT 5.330 931.545 1258.750 934.375 ;
        RECT 5.330 926.105 1258.750 928.935 ;
        RECT 5.330 920.665 1258.750 923.495 ;
        RECT 5.330 915.225 1258.750 918.055 ;
        RECT 5.330 909.785 1258.750 912.615 ;
        RECT 5.330 904.345 1258.750 907.175 ;
        RECT 5.330 898.905 1258.750 901.735 ;
        RECT 5.330 893.465 1258.750 896.295 ;
        RECT 5.330 888.025 1258.750 890.855 ;
        RECT 5.330 882.585 1258.750 885.415 ;
        RECT 5.330 877.145 1258.750 879.975 ;
        RECT 5.330 871.705 1258.750 874.535 ;
        RECT 5.330 866.265 1258.750 869.095 ;
        RECT 5.330 860.825 1258.750 863.655 ;
        RECT 5.330 855.385 1258.750 858.215 ;
        RECT 5.330 849.945 1258.750 852.775 ;
        RECT 5.330 844.505 1258.750 847.335 ;
        RECT 5.330 839.065 1258.750 841.895 ;
        RECT 5.330 833.625 1258.750 836.455 ;
        RECT 5.330 828.185 1258.750 831.015 ;
        RECT 5.330 822.745 1258.750 825.575 ;
        RECT 5.330 817.305 1258.750 820.135 ;
        RECT 5.330 811.865 1258.750 814.695 ;
        RECT 5.330 806.425 1258.750 809.255 ;
        RECT 5.330 800.985 1258.750 803.815 ;
        RECT 5.330 795.545 1258.750 798.375 ;
        RECT 5.330 790.105 1258.750 792.935 ;
        RECT 5.330 784.665 1258.750 787.495 ;
        RECT 5.330 779.225 1258.750 782.055 ;
        RECT 5.330 773.785 1258.750 776.615 ;
        RECT 5.330 768.345 1258.750 771.175 ;
        RECT 5.330 762.905 1258.750 765.735 ;
        RECT 5.330 757.465 1258.750 760.295 ;
        RECT 5.330 752.025 1258.750 754.855 ;
        RECT 5.330 746.585 1258.750 749.415 ;
        RECT 5.330 741.145 1258.750 743.975 ;
        RECT 5.330 735.705 1258.750 738.535 ;
        RECT 5.330 730.265 1258.750 733.095 ;
        RECT 5.330 724.825 1258.750 727.655 ;
        RECT 5.330 719.385 1258.750 722.215 ;
        RECT 5.330 713.945 1258.750 716.775 ;
        RECT 5.330 708.505 1258.750 711.335 ;
        RECT 5.330 703.065 1258.750 705.895 ;
        RECT 5.330 697.625 1258.750 700.455 ;
        RECT 5.330 692.185 1258.750 695.015 ;
        RECT 5.330 686.745 1258.750 689.575 ;
        RECT 5.330 681.305 1258.750 684.135 ;
        RECT 5.330 675.865 1258.750 678.695 ;
        RECT 5.330 670.425 1258.750 673.255 ;
        RECT 5.330 664.985 1258.750 667.815 ;
        RECT 5.330 659.545 1258.750 662.375 ;
        RECT 5.330 654.105 1258.750 656.935 ;
        RECT 5.330 648.665 1258.750 651.495 ;
        RECT 5.330 643.225 1258.750 646.055 ;
        RECT 5.330 637.785 1258.750 640.615 ;
        RECT 5.330 632.345 1258.750 635.175 ;
        RECT 5.330 626.905 1258.750 629.735 ;
        RECT 5.330 621.465 1258.750 624.295 ;
        RECT 5.330 616.025 1258.750 618.855 ;
        RECT 5.330 610.585 1258.750 613.415 ;
        RECT 5.330 605.145 1258.750 607.975 ;
        RECT 5.330 599.705 1258.750 602.535 ;
        RECT 5.330 594.265 1258.750 597.095 ;
        RECT 5.330 588.825 1258.750 591.655 ;
        RECT 5.330 583.385 1258.750 586.215 ;
        RECT 5.330 577.945 1258.750 580.775 ;
        RECT 5.330 572.505 1258.750 575.335 ;
        RECT 5.330 567.065 1258.750 569.895 ;
        RECT 5.330 561.625 1258.750 564.455 ;
        RECT 5.330 556.185 1258.750 559.015 ;
        RECT 5.330 550.745 1258.750 553.575 ;
        RECT 5.330 545.305 1258.750 548.135 ;
        RECT 5.330 539.865 1258.750 542.695 ;
        RECT 5.330 534.425 1258.750 537.255 ;
        RECT 5.330 528.985 1258.750 531.815 ;
        RECT 5.330 523.545 1258.750 526.375 ;
        RECT 5.330 518.105 1258.750 520.935 ;
        RECT 5.330 512.665 1258.750 515.495 ;
        RECT 5.330 507.225 1258.750 510.055 ;
        RECT 5.330 501.785 1258.750 504.615 ;
        RECT 5.330 496.345 1258.750 499.175 ;
        RECT 5.330 490.905 1258.750 493.735 ;
        RECT 5.330 485.465 1258.750 488.295 ;
        RECT 5.330 480.025 1258.750 482.855 ;
        RECT 5.330 474.585 1258.750 477.415 ;
        RECT 5.330 469.145 1258.750 471.975 ;
        RECT 5.330 463.705 1258.750 466.535 ;
        RECT 5.330 458.265 1258.750 461.095 ;
        RECT 5.330 452.825 1258.750 455.655 ;
        RECT 5.330 447.385 1258.750 450.215 ;
        RECT 5.330 441.945 1258.750 444.775 ;
        RECT 5.330 436.505 1258.750 439.335 ;
        RECT 5.330 431.065 1258.750 433.895 ;
        RECT 5.330 425.625 1258.750 428.455 ;
        RECT 5.330 420.185 1258.750 423.015 ;
        RECT 5.330 414.745 1258.750 417.575 ;
        RECT 5.330 409.305 1258.750 412.135 ;
        RECT 5.330 403.865 1258.750 406.695 ;
        RECT 5.330 398.425 1258.750 401.255 ;
        RECT 5.330 392.985 1258.750 395.815 ;
        RECT 5.330 387.545 1258.750 390.375 ;
        RECT 5.330 382.105 1258.750 384.935 ;
        RECT 5.330 376.665 1258.750 379.495 ;
        RECT 5.330 371.225 1258.750 374.055 ;
        RECT 5.330 365.785 1258.750 368.615 ;
        RECT 5.330 360.345 1258.750 363.175 ;
        RECT 5.330 354.905 1258.750 357.735 ;
        RECT 5.330 349.465 1258.750 352.295 ;
        RECT 5.330 344.025 1258.750 346.855 ;
        RECT 5.330 338.585 1258.750 341.415 ;
        RECT 5.330 333.145 1258.750 335.975 ;
        RECT 5.330 327.705 1258.750 330.535 ;
        RECT 5.330 322.265 1258.750 325.095 ;
        RECT 5.330 316.825 1258.750 319.655 ;
        RECT 5.330 311.385 1258.750 314.215 ;
        RECT 5.330 305.945 1258.750 308.775 ;
        RECT 5.330 300.505 1258.750 303.335 ;
        RECT 5.330 295.065 1258.750 297.895 ;
        RECT 5.330 289.625 1258.750 292.455 ;
        RECT 5.330 284.185 1258.750 287.015 ;
        RECT 5.330 278.745 1258.750 281.575 ;
        RECT 5.330 273.305 1258.750 276.135 ;
        RECT 5.330 267.865 1258.750 270.695 ;
        RECT 5.330 262.425 1258.750 265.255 ;
        RECT 5.330 256.985 1258.750 259.815 ;
        RECT 5.330 251.545 1258.750 254.375 ;
        RECT 5.330 246.105 1258.750 248.935 ;
        RECT 5.330 240.665 1258.750 243.495 ;
        RECT 5.330 235.225 1258.750 238.055 ;
        RECT 5.330 229.785 1258.750 232.615 ;
        RECT 5.330 224.345 1258.750 227.175 ;
        RECT 5.330 218.905 1258.750 221.735 ;
        RECT 5.330 213.465 1258.750 216.295 ;
        RECT 5.330 208.025 1258.750 210.855 ;
        RECT 5.330 202.585 1258.750 205.415 ;
        RECT 5.330 197.145 1258.750 199.975 ;
        RECT 5.330 191.705 1258.750 194.535 ;
        RECT 5.330 186.265 1258.750 189.095 ;
        RECT 5.330 180.825 1258.750 183.655 ;
        RECT 5.330 175.385 1258.750 178.215 ;
        RECT 5.330 169.945 1258.750 172.775 ;
        RECT 5.330 164.505 1258.750 167.335 ;
        RECT 5.330 159.065 1258.750 161.895 ;
        RECT 5.330 153.625 1258.750 156.455 ;
        RECT 5.330 148.185 1258.750 151.015 ;
        RECT 5.330 142.745 1258.750 145.575 ;
        RECT 5.330 137.305 1258.750 140.135 ;
        RECT 5.330 131.865 1258.750 134.695 ;
        RECT 5.330 126.425 1258.750 129.255 ;
        RECT 5.330 120.985 1258.750 123.815 ;
        RECT 5.330 115.545 1258.750 118.375 ;
        RECT 5.330 110.105 1258.750 112.935 ;
        RECT 5.330 104.665 1258.750 107.495 ;
        RECT 5.330 99.225 1258.750 102.055 ;
        RECT 5.330 93.785 1258.750 96.615 ;
        RECT 5.330 88.345 1258.750 91.175 ;
        RECT 5.330 82.905 1258.750 85.735 ;
        RECT 5.330 77.465 1258.750 80.295 ;
        RECT 5.330 72.025 1258.750 74.855 ;
        RECT 5.330 66.585 1258.750 69.415 ;
        RECT 5.330 61.145 1258.750 63.975 ;
        RECT 5.330 55.705 1258.750 58.535 ;
        RECT 5.330 50.265 1258.750 53.095 ;
        RECT 5.330 44.825 1258.750 47.655 ;
        RECT 5.330 39.385 1258.750 42.215 ;
        RECT 5.330 33.945 1258.750 36.775 ;
        RECT 5.330 28.505 1258.750 31.335 ;
        RECT 5.330 23.065 1258.750 25.895 ;
        RECT 5.330 17.625 1258.750 20.455 ;
        RECT 5.330 12.185 1258.750 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1258.560 1262.165 ;
      LAYER met1 ;
        RECT 5.520 5.480 1262.170 1262.320 ;
      LAYER met2 ;
        RECT 11.140 1270.880 315.830 1271.160 ;
        RECT 316.670 1270.880 947.870 1271.160 ;
        RECT 948.710 1270.880 1262.140 1271.160 ;
        RECT 11.140 4.280 1262.140 1270.880 ;
        RECT 11.140 3.670 27.870 4.280 ;
        RECT 28.710 3.670 39.370 4.280 ;
        RECT 40.210 3.670 50.870 4.280 ;
        RECT 51.710 3.670 62.370 4.280 ;
        RECT 63.210 3.670 73.870 4.280 ;
        RECT 74.710 3.670 85.370 4.280 ;
        RECT 86.210 3.670 96.870 4.280 ;
        RECT 97.710 3.670 108.370 4.280 ;
        RECT 109.210 3.670 119.870 4.280 ;
        RECT 120.710 3.670 131.370 4.280 ;
        RECT 132.210 3.670 142.870 4.280 ;
        RECT 143.710 3.670 154.370 4.280 ;
        RECT 155.210 3.670 165.870 4.280 ;
        RECT 166.710 3.670 177.370 4.280 ;
        RECT 178.210 3.670 188.870 4.280 ;
        RECT 189.710 3.670 200.370 4.280 ;
        RECT 201.210 3.670 211.870 4.280 ;
        RECT 212.710 3.670 223.370 4.280 ;
        RECT 224.210 3.670 234.870 4.280 ;
        RECT 235.710 3.670 246.370 4.280 ;
        RECT 247.210 3.670 257.870 4.280 ;
        RECT 258.710 3.670 269.370 4.280 ;
        RECT 270.210 3.670 280.870 4.280 ;
        RECT 281.710 3.670 292.370 4.280 ;
        RECT 293.210 3.670 303.870 4.280 ;
        RECT 304.710 3.670 315.370 4.280 ;
        RECT 316.210 3.670 326.870 4.280 ;
        RECT 327.710 3.670 338.370 4.280 ;
        RECT 339.210 3.670 349.870 4.280 ;
        RECT 350.710 3.670 361.370 4.280 ;
        RECT 362.210 3.670 372.870 4.280 ;
        RECT 373.710 3.670 384.370 4.280 ;
        RECT 385.210 3.670 395.870 4.280 ;
        RECT 396.710 3.670 407.370 4.280 ;
        RECT 408.210 3.670 418.870 4.280 ;
        RECT 419.710 3.670 430.370 4.280 ;
        RECT 431.210 3.670 441.870 4.280 ;
        RECT 442.710 3.670 453.370 4.280 ;
        RECT 454.210 3.670 464.870 4.280 ;
        RECT 465.710 3.670 476.370 4.280 ;
        RECT 477.210 3.670 487.870 4.280 ;
        RECT 488.710 3.670 499.370 4.280 ;
        RECT 500.210 3.670 510.870 4.280 ;
        RECT 511.710 3.670 522.370 4.280 ;
        RECT 523.210 3.670 533.870 4.280 ;
        RECT 534.710 3.670 545.370 4.280 ;
        RECT 546.210 3.670 556.870 4.280 ;
        RECT 557.710 3.670 568.370 4.280 ;
        RECT 569.210 3.670 579.870 4.280 ;
        RECT 580.710 3.670 591.370 4.280 ;
        RECT 592.210 3.670 602.870 4.280 ;
        RECT 603.710 3.670 614.370 4.280 ;
        RECT 615.210 3.670 625.870 4.280 ;
        RECT 626.710 3.670 637.370 4.280 ;
        RECT 638.210 3.670 648.870 4.280 ;
        RECT 649.710 3.670 660.370 4.280 ;
        RECT 661.210 3.670 671.870 4.280 ;
        RECT 672.710 3.670 683.370 4.280 ;
        RECT 684.210 3.670 694.870 4.280 ;
        RECT 695.710 3.670 706.370 4.280 ;
        RECT 707.210 3.670 717.870 4.280 ;
        RECT 718.710 3.670 729.370 4.280 ;
        RECT 730.210 3.670 740.870 4.280 ;
        RECT 741.710 3.670 752.370 4.280 ;
        RECT 753.210 3.670 763.870 4.280 ;
        RECT 764.710 3.670 775.370 4.280 ;
        RECT 776.210 3.670 786.870 4.280 ;
        RECT 787.710 3.670 798.370 4.280 ;
        RECT 799.210 3.670 809.870 4.280 ;
        RECT 810.710 3.670 821.370 4.280 ;
        RECT 822.210 3.670 832.870 4.280 ;
        RECT 833.710 3.670 844.370 4.280 ;
        RECT 845.210 3.670 855.870 4.280 ;
        RECT 856.710 3.670 867.370 4.280 ;
        RECT 868.210 3.670 878.870 4.280 ;
        RECT 879.710 3.670 890.370 4.280 ;
        RECT 891.210 3.670 901.870 4.280 ;
        RECT 902.710 3.670 913.370 4.280 ;
        RECT 914.210 3.670 924.870 4.280 ;
        RECT 925.710 3.670 936.370 4.280 ;
        RECT 937.210 3.670 947.870 4.280 ;
        RECT 948.710 3.670 959.370 4.280 ;
        RECT 960.210 3.670 970.870 4.280 ;
        RECT 971.710 3.670 982.370 4.280 ;
        RECT 983.210 3.670 993.870 4.280 ;
        RECT 994.710 3.670 1005.370 4.280 ;
        RECT 1006.210 3.670 1016.870 4.280 ;
        RECT 1017.710 3.670 1028.370 4.280 ;
        RECT 1029.210 3.670 1039.870 4.280 ;
        RECT 1040.710 3.670 1051.370 4.280 ;
        RECT 1052.210 3.670 1062.870 4.280 ;
        RECT 1063.710 3.670 1074.370 4.280 ;
        RECT 1075.210 3.670 1085.870 4.280 ;
        RECT 1086.710 3.670 1097.370 4.280 ;
        RECT 1098.210 3.670 1108.870 4.280 ;
        RECT 1109.710 3.670 1120.370 4.280 ;
        RECT 1121.210 3.670 1131.870 4.280 ;
        RECT 1132.710 3.670 1143.370 4.280 ;
        RECT 1144.210 3.670 1154.870 4.280 ;
        RECT 1155.710 3.670 1166.370 4.280 ;
        RECT 1167.210 3.670 1177.870 4.280 ;
        RECT 1178.710 3.670 1189.370 4.280 ;
        RECT 1190.210 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1212.370 4.280 ;
        RECT 1213.210 3.670 1223.870 4.280 ;
        RECT 1224.710 3.670 1235.370 4.280 ;
        RECT 1236.210 3.670 1262.140 4.280 ;
      LAYER met3 ;
        RECT 21.050 8.335 1253.895 1262.245 ;
      LAYER met4 ;
        RECT 25.135 19.895 97.440 1261.225 ;
        RECT 99.840 19.895 174.240 1261.225 ;
        RECT 176.640 19.895 251.040 1261.225 ;
        RECT 253.440 19.895 327.840 1261.225 ;
        RECT 330.240 19.895 404.640 1261.225 ;
        RECT 407.040 19.895 481.440 1261.225 ;
        RECT 483.840 19.895 558.240 1261.225 ;
        RECT 560.640 19.895 635.040 1261.225 ;
        RECT 637.440 19.895 711.840 1261.225 ;
        RECT 714.240 19.895 788.640 1261.225 ;
        RECT 791.040 19.895 865.440 1261.225 ;
        RECT 867.840 19.895 942.240 1261.225 ;
        RECT 944.640 19.895 1019.040 1261.225 ;
        RECT 1021.440 19.895 1095.840 1261.225 ;
        RECT 1098.240 19.895 1172.640 1261.225 ;
        RECT 1175.040 19.895 1249.440 1261.225 ;
        RECT 1251.840 19.895 1253.665 1261.225 ;
  END
END vco_adc_wrapper
END LIBRARY

