magic
tech sky130A
magscale 1 2
timestamp 1731453370
<< isosubstrate >>
rect 5100 -800 27000 -770
rect 4610 -1060 5020 -840
rect 5170 -1060 27000 -800
rect 4790 -5860 27000 -1060
rect 4790 -6000 5000 -5860
rect -10400 -6400 4490 -6000
rect 5330 -6040 27000 -5860
rect 5220 -6050 27000 -6040
rect 5020 -6400 27000 -6050
rect -10400 -24600 27000 -6400
<< locali >>
rect -710 8050 -310 8070
rect -710 8010 -690 8050
rect -650 8010 -610 8050
rect -570 8010 -530 8050
rect -490 8010 -450 8050
rect -410 8010 -370 8050
rect -330 8010 -310 8050
rect -710 7990 -310 8010
rect 3220 8050 3620 8070
rect 3220 8010 3240 8050
rect 3280 8010 3320 8050
rect 3360 8010 3400 8050
rect 3440 8010 3480 8050
rect 3520 8010 3560 8050
rect 3600 8010 3620 8050
rect 3220 7990 3620 8010
rect -2800 4070 -1030 4090
rect -2800 4030 -1210 4070
rect -1170 4030 -1130 4070
rect -1090 4030 -1030 4070
rect -2800 3990 -2780 4030
rect -2740 3990 -2700 4030
rect -2660 3990 -1030 4030
rect -2800 3950 -1210 3990
rect -1170 3950 -1130 3990
rect -1090 3950 -1030 3990
rect -2800 3910 -2780 3950
rect -2740 3910 -2700 3950
rect -2660 3910 -1030 3950
rect -2800 3890 -1030 3910
rect 1850 4070 2050 4090
rect 1850 4010 1870 4070
rect 1930 4010 1970 4070
rect 2030 4010 2050 4070
rect 1850 3970 2050 4010
rect 1850 3910 1870 3970
rect 1930 3910 1970 3970
rect 2030 3910 2050 3970
rect 2870 4010 3050 4030
rect 2870 3960 2880 4010
rect 2930 3960 2980 4010
rect 3030 3960 3050 4010
rect 2870 3930 3050 3960
rect 1850 3890 2050 3910
rect 1890 1570 2000 3890
rect 1890 1510 1920 1570
rect 1980 1510 2000 1570
rect 1890 1450 2000 1510
rect 1890 1390 1920 1450
rect 1980 1390 2000 1450
rect 1890 1370 2000 1390
rect 5980 -1160 6100 -1140
rect 5980 -1210 6000 -1160
rect 6050 -1210 6100 -1160
rect 5980 -1230 6100 -1210
rect 5980 -1260 7180 -1230
rect 5980 -1310 6000 -1260
rect 6050 -1310 6100 -1260
rect 6150 -1310 7180 -1260
rect 5980 -1330 7180 -1310
rect 1130 -1560 6110 -1540
rect 1130 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 1130 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 6030 -1700 6110 -1680
rect 7080 -1650 7180 -1330
rect 7080 -1680 7320 -1650
rect 7080 -1720 7100 -1680
rect 7140 -1720 7180 -1680
rect 7220 -1720 7260 -1680
rect 7300 -1720 7320 -1680
rect 7080 -1760 7320 -1720
rect 1470 -2150 2740 -2130
rect 1470 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 1470 -2220 2740 -2210
rect 1530 -2230 2740 -2220
rect 1580 -2410 4120 -2380
rect 1580 -2470 3910 -2410
rect 3970 -2470 4030 -2410
rect 4090 -2470 4120 -2410
rect 1580 -2500 4120 -2470
rect 4000 -2530 4120 -2500
rect 4000 -2590 4030 -2530
rect 4090 -2590 4120 -2530
rect 4000 -2620 4120 -2590
rect 4000 -4770 4120 -4740
rect 4000 -4830 4030 -4770
rect 4090 -4830 4120 -4770
rect 4000 -4860 4120 -4830
rect 2060 -4890 4120 -4860
rect 2060 -4950 2080 -4890
rect 2140 -4950 2200 -4890
rect 2260 -4950 2320 -4890
rect 2380 -4950 3900 -4890
rect 3960 -4950 4030 -4890
rect 4090 -4950 4120 -4890
rect 2060 -4980 4120 -4950
rect 4000 -5010 4120 -4980
rect 850 -6110 1050 -5060
rect 4000 -5070 4030 -5010
rect 4090 -5070 4120 -5010
rect 4000 -5100 4120 -5070
rect 850 -6190 3280 -6110
rect 850 -6250 2910 -6190
rect 2970 -6250 3030 -6190
rect 3090 -6250 3150 -6190
rect 3210 -6250 3280 -6190
rect 850 -6310 3280 -6250
rect -2240 -6750 -1830 -6740
rect -2240 -6760 -1820 -6750
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -1820 -6760
rect -2240 -6820 -1820 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -2240 -6900 -2160 -6880
rect -2800 -7800 -1860 -7780
rect -2800 -7840 -2780 -7800
rect -2740 -7840 -2700 -7800
rect -2660 -7840 -2620 -7800
rect -2580 -7840 -2080 -7800
rect -2040 -7840 -2000 -7800
rect -1960 -7840 -1920 -7800
rect -1880 -7840 -1860 -7800
rect -2800 -7860 -1860 -7840
rect 1260 -7890 2370 -7870
rect 1260 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 1260 -7950 2370 -7930
rect 16510 -7970 16600 -7870
rect 16650 -7900 17170 -7870
rect 16650 -7940 16680 -7900
rect 16720 -7940 17170 -7900
rect 16650 -7970 17170 -7940
rect 4000 -8620 4120 -8590
rect 4000 -8680 4030 -8620
rect 4090 -8680 4120 -8620
rect 4000 -8710 4120 -8680
rect 1580 -8740 4120 -8710
rect 1580 -8800 3900 -8740
rect 3960 -8800 4030 -8740
rect 4090 -8800 4120 -8740
rect 1580 -8830 4120 -8800
rect -1640 -9140 -1380 -9100
rect -2400 -9360 -1380 -9140
rect -2400 -9380 -1800 -9360
rect -1840 -9420 -1800 -9380
rect -1740 -9420 -1680 -9360
rect -1620 -9420 -1380 -9360
rect -1840 -9480 -1380 -9420
rect -1840 -9540 -1800 -9480
rect -1740 -9540 -1680 -9480
rect -1620 -9540 -1380 -9480
rect -1840 -9560 -1380 -9540
rect 17070 -9960 17170 -7970
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect 17000 -10040 17170 -10020
rect 17000 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect 17000 -10100 17170 -10080
<< viali >>
rect -690 8010 -650 8050
rect -610 8010 -570 8050
rect -530 8010 -490 8050
rect -450 8010 -410 8050
rect -370 8010 -330 8050
rect 3240 8010 3280 8050
rect 3320 8010 3360 8050
rect 3400 8010 3440 8050
rect 3480 8010 3520 8050
rect 3560 8010 3600 8050
rect 11060 8010 11100 8050
rect 11140 8010 11180 8050
rect 11220 8010 11260 8050
rect 11300 8010 11340 8050
rect 11380 8010 11420 8050
rect 15890 8010 15930 8050
rect 15970 8010 16010 8050
rect 16050 8010 16090 8050
rect 16130 8010 16170 8050
rect 16210 8010 16250 8050
rect -1210 4030 -1170 4070
rect -1130 4030 -1090 4070
rect -2780 3990 -2740 4030
rect -2700 3990 -2660 4030
rect -1210 3950 -1170 3990
rect -1130 3950 -1090 3990
rect -2780 3910 -2740 3950
rect -2700 3910 -2660 3950
rect 1870 4010 1930 4070
rect 1970 4010 2030 4070
rect 1870 3910 1930 3970
rect 1970 3910 2030 3970
rect 2880 3960 2930 4010
rect 2980 3960 3030 4010
rect 1920 1510 1980 1570
rect 1920 1390 1980 1450
rect -2000 -470 -1960 -430
rect -1920 -470 -1880 -430
rect 6000 -1210 6050 -1160
rect 6000 -1310 6050 -1260
rect 6100 -1310 6150 -1260
rect 1150 -1600 1190 -1560
rect 1230 -1600 1270 -1560
rect 5970 -1600 6010 -1560
rect 6050 -1600 6090 -1560
rect 6050 -1680 6090 -1640
rect 7100 -1720 7140 -1680
rect 7180 -1720 7220 -1680
rect 7260 -1720 7300 -1680
rect 2420 -2210 2480 -2150
rect 2540 -2210 2600 -2150
rect 2660 -2210 2720 -2150
rect 3910 -2470 3970 -2410
rect 4030 -2470 4090 -2410
rect 4030 -2590 4090 -2530
rect 4030 -4830 4090 -4770
rect 2080 -4950 2140 -4890
rect 2200 -4950 2260 -4890
rect 2320 -4950 2380 -4890
rect 3900 -4950 3960 -4890
rect 4030 -4950 4090 -4890
rect 4030 -5070 4090 -5010
rect 2910 -6250 2970 -6190
rect 3030 -6250 3090 -6190
rect 3150 -6250 3210 -6190
rect -2220 -6800 -2180 -6760
rect -2140 -6800 -2100 -6760
rect -2220 -6880 -2180 -6840
rect -2780 -7840 -2740 -7800
rect -2700 -7840 -2660 -7800
rect -2620 -7840 -2580 -7800
rect -2080 -7840 -2040 -7800
rect -2000 -7840 -1960 -7800
rect -1920 -7840 -1880 -7800
rect 1280 -7930 1320 -7890
rect 1360 -7930 1400 -7890
rect 1440 -7930 1480 -7890
rect 2150 -7930 2190 -7890
rect 2230 -7930 2270 -7890
rect 2310 -7930 2350 -7890
rect 16680 -7940 16720 -7900
rect 4030 -8680 4090 -8620
rect 3900 -8800 3960 -8740
rect 4030 -8800 4090 -8740
rect -1800 -9420 -1740 -9360
rect -1680 -9420 -1620 -9360
rect -1800 -9540 -1740 -9480
rect -1680 -9540 -1620 -9480
rect 17100 -10000 17140 -9960
rect 17020 -10080 17060 -10040
rect 17100 -10080 17140 -10040
<< metal1 >>
rect -710 8060 -310 8070
rect -710 8000 -700 8060
rect -640 8050 -580 8060
rect -520 8050 -460 8060
rect -400 8050 -310 8060
rect -640 8010 -610 8050
rect -490 8010 -460 8050
rect -400 8010 -370 8050
rect -330 8010 -310 8050
rect -640 8000 -580 8010
rect -520 8000 -460 8010
rect -400 8000 -310 8010
rect -710 7990 -310 8000
rect 3220 8060 3620 8070
rect 3220 8000 3230 8060
rect 3290 8050 3390 8060
rect 3450 8050 3550 8060
rect 3290 8010 3320 8050
rect 3360 8010 3390 8050
rect 3450 8010 3480 8050
rect 3520 8010 3550 8050
rect 3290 8000 3390 8010
rect 3450 8000 3550 8010
rect 3610 8000 3620 8060
rect 3220 7990 3620 8000
rect 11040 8060 11440 8070
rect 11040 8000 11050 8060
rect 11110 8050 11210 8060
rect 11270 8050 11370 8060
rect 11110 8010 11140 8050
rect 11180 8010 11210 8050
rect 11270 8010 11300 8050
rect 11340 8010 11370 8050
rect 11110 8000 11210 8010
rect 11270 8000 11370 8010
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8060 16270 8070
rect 15870 8000 15880 8060
rect 15940 8050 16040 8060
rect 16100 8050 16200 8060
rect 15940 8010 15970 8050
rect 16010 8010 16040 8050
rect 16100 8010 16130 8050
rect 16170 8010 16200 8050
rect 15940 8000 16040 8010
rect 16100 8000 16200 8010
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 6890 4900 7140 4960
rect 6890 4840 6910 4900
rect 6970 4840 7030 4900
rect 7090 4840 7140 4900
rect 6890 4800 7140 4840
rect -2800 4030 -2600 4090
rect -2800 3990 -2780 4030
rect -2740 3990 -2700 4030
rect -2660 3990 -2600 4030
rect -2800 3950 -2600 3990
rect -2800 3910 -2780 3950
rect -2740 3910 -2700 3950
rect -2660 3910 -2600 3950
rect -2800 -1450 -2600 3910
rect -1230 4070 3050 4090
rect -1230 4030 -1210 4070
rect -1170 4030 -1130 4070
rect -1090 4030 1870 4070
rect -1230 4010 1870 4030
rect 1930 4010 1970 4070
rect 2030 4010 3050 4070
rect -1230 3990 2880 4010
rect -1230 3950 -1210 3990
rect -1170 3950 -1130 3990
rect -1090 3970 2880 3990
rect -1090 3950 1870 3970
rect -1230 3910 1870 3950
rect 1930 3910 1970 3970
rect 2030 3960 2880 3970
rect 2930 3960 2980 4010
rect 3030 3960 3050 4010
rect 2030 3910 3050 3960
rect -1230 3890 3050 3910
rect -2020 -410 -1920 2100
rect 1890 1570 2000 1590
rect 1890 1510 1920 1570
rect 1980 1510 2000 1570
rect 1890 1450 2000 1510
rect 1890 1390 1920 1450
rect 1980 1390 2000 1450
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 -130 -1080 1010
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 -120 80 1000
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 -130 1290 1020
rect 1890 1030 2000 1390
rect 1890 910 6100 1030
rect -2020 -430 -1860 -410
rect -2020 -470 -2000 -430
rect -1960 -470 -1920 -430
rect -1880 -470 -1860 -430
rect -2020 -490 -1860 -470
rect 5980 -1160 6100 910
rect 5980 -1210 6000 -1160
rect 6050 -1210 6100 -1160
rect 5980 -1230 6100 -1210
rect 5980 -1260 6170 -1230
rect 5980 -1310 6000 -1260
rect 6050 -1310 6100 -1260
rect 6150 -1310 6170 -1260
rect 5980 -1330 6170 -1310
rect -2800 -1530 -1720 -1450
rect -2800 -7780 -2600 -1530
rect 970 -1560 1290 -1540
rect 970 -1600 1150 -1560
rect 1190 -1600 1230 -1560
rect 1270 -1600 1290 -1560
rect 970 -1620 1290 -1600
rect 5950 -1560 6110 -1540
rect 5950 -1600 5970 -1560
rect 6010 -1600 6050 -1560
rect 6090 -1600 6110 -1560
rect 5950 -1620 6110 -1600
rect 6030 -1640 6110 -1620
rect 6030 -1680 6050 -1640
rect 6090 -1680 6110 -1640
rect 2400 -2150 2740 -2130
rect 2400 -2210 2420 -2150
rect 2480 -2210 2540 -2150
rect 2600 -2210 2660 -2150
rect 2720 -2210 2740 -2150
rect 2400 -2230 2740 -2210
rect 2360 -3100 2760 -2230
rect 3880 -2410 4120 -2380
rect 3880 -2470 3910 -2410
rect 3970 -2470 4030 -2410
rect 4090 -2470 4120 -2410
rect 3880 -2500 4120 -2470
rect 4000 -2530 4120 -2500
rect 4000 -2590 4030 -2530
rect 4090 -2590 4120 -2530
rect 4000 -2730 4120 -2590
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3480 2760 -3280
rect -2320 -4490 -1920 -3900
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4800 -1920 -4550
rect -1770 -4210 -1570 -4190
rect -1770 -4270 -1710 -4210
rect -1650 -4270 -1570 -4210
rect -1770 -4330 -1570 -4270
rect -1770 -4390 -1710 -4330
rect -1650 -4390 -1570 -4330
rect -1770 -4450 -1570 -4390
rect -1770 -4510 -1710 -4450
rect -1650 -4510 -1570 -4450
rect -1770 -4570 -1570 -4510
rect -1770 -4630 -1710 -4570
rect -1650 -4630 -1570 -4570
rect -1770 -4660 -1570 -4630
rect 4001 -4740 4120 -2730
rect 4000 -4770 4120 -4740
rect 4000 -4830 4030 -4770
rect 4090 -4830 4120 -4770
rect 4000 -4860 4120 -4830
rect 2060 -4890 2420 -4860
rect 2060 -4950 2080 -4890
rect 2140 -4950 2200 -4890
rect 2260 -4950 2320 -4890
rect 2380 -4950 2420 -4890
rect 2060 -4980 2420 -4950
rect 3880 -4890 4120 -4860
rect 3880 -4950 3900 -4890
rect 3960 -4950 4030 -4890
rect 4090 -4950 4120 -4890
rect 6030 -4830 6110 -1680
rect 7080 -1680 8560 -1650
rect 7080 -1720 7100 -1680
rect 7140 -1720 7180 -1680
rect 7220 -1720 7260 -1680
rect 7300 -1720 8560 -1680
rect 7080 -1760 8560 -1720
rect 18510 -2410 18610 -2340
rect 18510 -2470 18530 -2410
rect 18590 -2470 18610 -2410
rect 18510 -2530 18610 -2470
rect 18510 -2590 18530 -2530
rect 18590 -2590 18610 -2530
rect 18510 -2650 18610 -2590
rect 18510 -2710 18530 -2650
rect 18590 -2710 18610 -2650
rect 18510 -2740 18610 -2710
rect 13160 -3580 13250 -3540
rect 13160 -3640 13170 -3580
rect 13230 -3640 13250 -3580
rect 13160 -3700 13250 -3640
rect 13160 -3760 13170 -3700
rect 13230 -3760 13250 -3700
rect 13160 -3890 13250 -3760
rect 7000 -4420 7220 -4400
rect 7000 -4480 7020 -4420
rect 7080 -4480 7140 -4420
rect 7200 -4480 7220 -4420
rect 7000 -4500 7220 -4480
rect 7000 -4540 8240 -4500
rect 7000 -4600 7020 -4540
rect 7080 -4600 7140 -4540
rect 7200 -4600 8240 -4540
rect 7000 -4620 7220 -4600
rect 6030 -4910 6520 -4830
rect 3880 -4980 4120 -4950
rect 4000 -5010 4120 -4980
rect -1790 -6070 -1710 -5020
rect 4000 -5070 4030 -5010
rect 4090 -5070 4120 -5010
rect 4000 -5100 4120 -5070
rect -1480 -5500 -1080 -5340
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5580 -1080 -5560
rect 250 -5500 650 -5330
rect 250 -5560 280 -5500
rect 340 -5560 400 -5500
rect 460 -5560 520 -5500
rect 580 -5560 650 -5500
rect 250 -5580 650 -5560
rect 2090 -5500 2490 -5330
rect 2090 -5560 2120 -5500
rect 2180 -5560 2240 -5500
rect 2300 -5560 2360 -5500
rect 2420 -5560 2490 -5500
rect 2090 -5580 2490 -5560
rect -1790 -6150 2370 -6070
rect -2240 -6760 -2080 -6740
rect -2240 -6800 -2220 -6760
rect -2180 -6800 -2140 -6760
rect -2100 -6800 -2080 -6760
rect -2240 -6820 -2080 -6800
rect -2240 -6840 -2160 -6820
rect -2240 -6880 -2220 -6840
rect -2180 -6880 -2160 -6840
rect -2800 -7800 -2560 -7780
rect -2800 -7840 -2780 -7800
rect -2740 -7840 -2700 -7800
rect -2660 -7840 -2620 -7800
rect -2580 -7840 -2560 -7800
rect -2800 -7860 -2560 -7840
rect -2800 -7910 -2600 -7860
rect -2800 -7970 -2730 -7910
rect -2670 -7970 -2600 -7910
rect -2800 -8030 -2600 -7970
rect -2800 -8090 -2730 -8030
rect -2670 -8090 -2600 -8030
rect -2800 -8150 -2600 -8090
rect -2800 -8210 -2730 -8150
rect -2670 -8210 -2600 -8150
rect -2800 -8240 -2600 -8210
rect -2240 -10020 -2160 -6880
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7170 -1480 -7150
rect -2100 -7800 -1720 -7780
rect -2100 -7840 -2080 -7800
rect -2040 -7840 -2000 -7800
rect -1960 -7840 -1920 -7800
rect -1880 -7840 -1720 -7800
rect -2100 -7860 -1720 -7840
rect 2290 -7870 2370 -6150
rect 2880 -6190 3280 -6110
rect 2880 -6250 2910 -6190
rect 2970 -6250 3030 -6190
rect 3090 -6250 3150 -6190
rect 3210 -6250 3280 -6190
rect 2880 -6360 3280 -6250
rect 2880 -6460 2920 -6360
rect 3020 -6460 3120 -6360
rect 3220 -6460 3280 -6360
rect 2880 -6530 3280 -6460
rect 2880 -6630 3020 -6530
rect 3120 -6630 3280 -6530
rect 2880 -6690 3280 -6630
rect 970 -7890 1500 -7870
rect 970 -7930 1280 -7890
rect 1320 -7930 1360 -7890
rect 1400 -7930 1440 -7890
rect 1480 -7930 1500 -7890
rect 970 -7950 1500 -7930
rect 2130 -7890 2370 -7870
rect 2130 -7930 2150 -7890
rect 2190 -7930 2230 -7890
rect 2270 -7930 2310 -7890
rect 2350 -7930 2370 -7890
rect 2130 -7950 2370 -7930
rect 4001 -8590 4120 -5100
rect 6440 -7010 6520 -4910
rect 9110 -4950 9310 -4930
rect 9110 -5010 9130 -4950
rect 9190 -5010 9230 -4950
rect 9290 -5010 9310 -4950
rect 9110 -5050 9310 -5010
rect 9110 -5110 9130 -5050
rect 9190 -5110 9230 -5050
rect 9290 -5110 9310 -5050
rect 9110 -5130 9310 -5110
rect 16280 -7900 16750 -7870
rect 16280 -7940 16680 -7900
rect 16720 -7940 16750 -7900
rect 16280 -7970 16750 -7940
rect 4000 -8620 4120 -8590
rect 4000 -8680 4030 -8620
rect 4090 -8680 4120 -8620
rect 4000 -8710 4120 -8680
rect 3880 -8740 4120 -8710
rect 3880 -8800 3900 -8740
rect 3960 -8800 4030 -8740
rect 4090 -8800 4120 -8740
rect 3880 -8830 4120 -8800
rect -1640 -9140 -1240 -9050
rect 580 -9140 980 -9060
rect -150 -9160 250 -9140
rect -150 -9220 -120 -9160
rect -60 -9220 0 -9160
rect 60 -9220 120 -9160
rect 180 -9220 250 -9160
rect -150 -9250 250 -9220
rect -1840 -9360 -1600 -9320
rect -1840 -9420 -1800 -9360
rect -1740 -9420 -1680 -9360
rect -1620 -9420 -1600 -9360
rect -1840 -9480 -1600 -9420
rect -1840 -9540 -1800 -9480
rect -1740 -9540 -1680 -9480
rect -1620 -9540 -1600 -9480
rect -1840 -9570 -1440 -9540
rect -1840 -9630 -1810 -9570
rect -1750 -9630 -1690 -9570
rect -1630 -9630 -1570 -9570
rect -1510 -9630 -1440 -9570
rect -1840 -9770 -1440 -9630
rect 17070 -9960 17170 -9940
rect 17070 -10000 17100 -9960
rect 17140 -10000 17170 -9960
rect 17070 -10020 17170 -10000
rect -2240 -10040 17170 -10020
rect -2240 -10080 17020 -10040
rect 17060 -10080 17100 -10040
rect 17140 -10080 17170 -10040
rect -2240 -10100 17170 -10080
<< via1 >>
rect -700 8050 -640 8060
rect -580 8050 -520 8060
rect -460 8050 -400 8060
rect -700 8010 -690 8050
rect -690 8010 -650 8050
rect -650 8010 -640 8050
rect -580 8010 -570 8050
rect -570 8010 -530 8050
rect -530 8010 -520 8050
rect -460 8010 -450 8050
rect -450 8010 -410 8050
rect -410 8010 -400 8050
rect -700 8000 -640 8010
rect -580 8000 -520 8010
rect -460 8000 -400 8010
rect 3230 8050 3290 8060
rect 3390 8050 3450 8060
rect 3550 8050 3610 8060
rect 3230 8010 3240 8050
rect 3240 8010 3280 8050
rect 3280 8010 3290 8050
rect 3390 8010 3400 8050
rect 3400 8010 3440 8050
rect 3440 8010 3450 8050
rect 3550 8010 3560 8050
rect 3560 8010 3600 8050
rect 3600 8010 3610 8050
rect 3230 8000 3290 8010
rect 3390 8000 3450 8010
rect 3550 8000 3610 8010
rect 11050 8050 11110 8060
rect 11210 8050 11270 8060
rect 11370 8050 11430 8060
rect 11050 8010 11060 8050
rect 11060 8010 11100 8050
rect 11100 8010 11110 8050
rect 11210 8010 11220 8050
rect 11220 8010 11260 8050
rect 11260 8010 11270 8050
rect 11370 8010 11380 8050
rect 11380 8010 11420 8050
rect 11420 8010 11430 8050
rect 11050 8000 11110 8010
rect 11210 8000 11270 8010
rect 11370 8000 11430 8010
rect 15880 8050 15940 8060
rect 16040 8050 16100 8060
rect 16200 8050 16260 8060
rect 15880 8010 15890 8050
rect 15890 8010 15930 8050
rect 15930 8010 15940 8050
rect 16040 8010 16050 8050
rect 16050 8010 16090 8050
rect 16090 8010 16100 8050
rect 16200 8010 16210 8050
rect 16210 8010 16250 8050
rect 16250 8010 16260 8050
rect 15880 8000 15940 8010
rect 16040 8000 16100 8010
rect 16200 8000 16260 8010
rect 6910 4840 6970 4900
rect 7030 4840 7090 4900
rect 14700 4570 14760 4630
rect 14700 4450 14760 4510
rect 14700 4330 14760 4390
rect -1430 1010 -1360 1080
rect -1200 1010 -1130 1080
rect -270 1000 -200 1070
rect -50 1000 20 1070
rect 930 1020 990 1080
rect 1180 1020 1240 1080
rect 2390 -3160 2450 -3100
rect 2510 -3160 2570 -3100
rect 2630 -3160 2690 -3100
rect 2390 -3280 2450 -3220
rect 2510 -3280 2570 -3220
rect 2630 -3280 2690 -3220
rect -2280 -4550 -2220 -4490
rect -2030 -4550 -1970 -4490
rect -1710 -4270 -1650 -4210
rect -1710 -4390 -1650 -4330
rect -1710 -4510 -1650 -4450
rect -1710 -4630 -1650 -4570
rect 18530 -2470 18590 -2410
rect 18530 -2590 18590 -2530
rect 18530 -2710 18590 -2650
rect 13170 -3640 13230 -3580
rect 13170 -3760 13230 -3700
rect 7020 -4480 7080 -4420
rect 7140 -4480 7200 -4420
rect 7020 -4600 7080 -4540
rect 7140 -4600 7200 -4540
rect -1450 -5560 -1390 -5500
rect -1330 -5560 -1270 -5500
rect -1210 -5560 -1150 -5500
rect 280 -5560 340 -5500
rect 400 -5560 460 -5500
rect 520 -5560 580 -5500
rect 2120 -5560 2180 -5500
rect 2240 -5560 2300 -5500
rect 2360 -5560 2420 -5500
rect -2730 -7970 -2670 -7910
rect -2730 -8090 -2670 -8030
rect -2730 -8210 -2670 -8150
rect -1930 -7150 -1870 -7090
rect -1810 -7150 -1750 -7090
rect -1690 -7150 -1630 -7090
rect -1570 -7150 -1510 -7090
rect 2920 -6460 3020 -6360
rect 3120 -6460 3220 -6360
rect 3020 -6630 3120 -6530
rect 9130 -5010 9190 -4950
rect 9230 -5010 9290 -4950
rect 9130 -5110 9190 -5050
rect 9230 -5110 9290 -5050
rect 18530 -7070 18590 -7010
rect 18530 -7190 18590 -7130
rect 18530 -7310 18590 -7250
rect -120 -9220 -60 -9160
rect 0 -9220 60 -9160
rect 120 -9220 180 -9160
rect -1810 -9630 -1750 -9570
rect -1690 -9630 -1630 -9570
rect -1570 -9630 -1510 -9570
rect 10030 -9640 10090 -9580
rect 10150 -9640 10210 -9580
rect 10270 -9640 10330 -9580
rect 16090 -9640 16150 -9580
rect 16210 -9640 16270 -9580
rect 16330 -9640 16390 -9580
<< metal2 >>
rect 39514 32062 41630 32430
rect -710 8180 -310 8210
rect -710 8100 -670 8180
rect -590 8100 -430 8180
rect -350 8100 -310 8180
rect -710 8060 -310 8100
rect -710 8000 -700 8060
rect -640 8000 -580 8060
rect -520 8000 -460 8060
rect -400 8000 -310 8060
rect -710 7990 -310 8000
rect 3220 8190 3620 8210
rect 3220 8110 3260 8190
rect 3340 8110 3480 8190
rect 3560 8110 3620 8190
rect 3220 8060 3620 8110
rect 3220 8000 3230 8060
rect 3290 8000 3390 8060
rect 3450 8000 3550 8060
rect 3610 8000 3620 8060
rect 3220 7990 3620 8000
rect 11040 8190 11440 8220
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8060 11440 8110
rect 11040 8000 11050 8060
rect 11110 8000 11210 8060
rect 11270 8000 11370 8060
rect 11430 8000 11440 8060
rect 11040 7990 11440 8000
rect 15870 8180 16270 8210
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8060 16270 8100
rect 15870 8000 15880 8060
rect 15940 8000 16040 8060
rect 16100 8000 16200 8060
rect 16260 8000 16270 8060
rect 15870 7990 16270 8000
rect 39490 5100 39890 32062
rect 20600 5000 39890 5100
rect 7140 4960 39890 5000
rect 6890 4900 39890 4960
rect 6890 4840 6910 4900
rect 6970 4840 7030 4900
rect 7090 4840 39890 4900
rect 6890 4800 39890 4840
rect 20600 4700 39890 4800
rect 14680 4640 14990 4700
rect 14680 4630 14830 4640
rect 14680 4570 14700 4630
rect 14760 4570 14830 4630
rect 14680 4540 14830 4570
rect 14930 4540 14990 4640
rect 14680 4510 14990 4540
rect 14680 4450 14700 4510
rect 14760 4450 14990 4510
rect 14680 4440 14990 4450
rect 14680 4390 14830 4440
rect 14680 4330 14700 4390
rect 14760 4340 14830 4390
rect 14930 4340 14990 4440
rect 14760 4330 14990 4340
rect 14680 4300 14990 4330
rect -1480 1080 -1080 1110
rect -1480 1010 -1430 1080
rect -1360 1010 -1200 1080
rect -1130 1010 -1080 1080
rect -1480 960 -1080 1010
rect -1480 880 -1430 960
rect -1350 880 -1220 960
rect -1140 880 -1080 960
rect -1480 820 -1080 880
rect -1480 740 -1430 820
rect -1350 740 -1220 820
rect -1140 740 -1080 820
rect -1480 710 -1080 740
rect -320 1070 80 1110
rect -320 1000 -270 1070
rect -200 1000 -50 1070
rect 20 1000 80 1070
rect -320 950 80 1000
rect -320 870 -270 950
rect -190 870 -50 950
rect 30 870 80 950
rect -320 810 80 870
rect -320 730 -270 810
rect -190 730 -50 810
rect 30 730 80 810
rect -320 710 80 730
rect 890 1080 1290 1110
rect 890 1020 930 1080
rect 990 1020 1180 1080
rect 1240 1020 1290 1080
rect 890 980 1290 1020
rect 890 900 930 980
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 890 820 1290 900
rect 890 740 930 820
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 890 710 1290 740
rect 4610 -900 5020 -840
rect 4610 -1000 4650 -900
rect 4750 -1000 4860 -900
rect 4960 -1000 5020 -900
rect 4610 -1060 5020 -1000
rect 4800 -1110 5020 -1060
rect 4800 -1210 4860 -1110
rect 4960 -1210 5020 -1110
rect 2360 -3100 2760 -3080
rect 2360 -3160 2390 -3100
rect 2450 -3160 2510 -3100
rect 2570 -3160 2630 -3100
rect 2690 -3160 2760 -3100
rect 2360 -3220 2760 -3160
rect 2360 -3280 2390 -3220
rect 2450 -3280 2510 -3220
rect 2570 -3280 2630 -3220
rect 2690 -3280 2760 -3220
rect 2360 -3340 2760 -3280
rect 2360 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect 2360 -3430 2760 -3420
rect -2320 -4220 -1920 -4190
rect -2320 -4300 -2290 -4220
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -2320 -4370 -1920 -4300
rect -2320 -4450 -2290 -4370
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -2320 -4490 -1920 -4450
rect -2320 -4550 -2280 -4490
rect -2220 -4550 -2030 -4490
rect -1970 -4550 -1920 -4490
rect -2320 -4590 -1920 -4550
rect -1770 -4210 -1570 -4190
rect -1770 -4270 -1710 -4210
rect -1650 -4270 -1570 -4210
rect -1770 -4330 -1570 -4270
rect -1770 -4390 -1710 -4330
rect -1650 -4390 -1570 -4330
rect -1770 -4450 -1570 -4390
rect -1770 -4510 -1710 -4450
rect -1650 -4510 -1570 -4450
rect -1770 -4570 -1570 -4510
rect -1770 -4630 -1710 -4570
rect -1650 -4630 -1570 -4570
rect 4800 -4400 5020 -1210
rect 18510 -2390 18790 -2340
rect 18510 -2410 18650 -2390
rect 18510 -2470 18530 -2410
rect 18590 -2470 18650 -2410
rect 18730 -2470 18790 -2390
rect 18510 -2530 18790 -2470
rect 18510 -2590 18530 -2530
rect 18590 -2550 18790 -2530
rect 18590 -2590 18650 -2550
rect 18510 -2630 18650 -2590
rect 18730 -2630 18790 -2550
rect 18510 -2650 18790 -2630
rect 18510 -2710 18530 -2650
rect 18590 -2710 18790 -2650
rect 18510 -2740 18790 -2710
rect 13160 -3570 13420 -3540
rect 13160 -3580 13300 -3570
rect 13160 -3640 13170 -3580
rect 13230 -3640 13300 -3580
rect 13160 -3650 13300 -3640
rect 13380 -3650 13420 -3570
rect 13160 -3700 13420 -3650
rect 13160 -3760 13170 -3700
rect 13230 -3760 13420 -3700
rect 13160 -3810 13420 -3760
rect 13160 -3890 13300 -3810
rect 13380 -3890 13420 -3810
rect 13160 -3940 13420 -3890
rect 4800 -4420 7220 -4400
rect 4800 -4480 7020 -4420
rect 7080 -4480 7140 -4420
rect 7200 -4480 7220 -4420
rect 4800 -4540 7220 -4480
rect 4800 -4600 7020 -4540
rect 7080 -4600 7140 -4540
rect 7200 -4600 7220 -4540
rect 4800 -4620 7220 -4600
rect -1770 -4800 -1570 -4630
rect -7380 -5000 -1570 -4800
rect 9110 -4950 9310 -4930
rect -7380 -25254 -6980 -5000
rect 9110 -5010 9130 -4950
rect 9190 -5010 9230 -4950
rect 9290 -5010 9310 -4950
rect 9110 -5050 9310 -5010
rect 9110 -5110 9130 -5050
rect 9190 -5110 9230 -5050
rect 9290 -5110 9310 -5050
rect -1480 -5500 -1080 -5470
rect -1480 -5560 -1450 -5500
rect -1390 -5560 -1330 -5500
rect -1270 -5560 -1210 -5500
rect -1150 -5560 -1080 -5500
rect -1480 -5630 -1080 -5560
rect -1480 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 -1080 -5630
rect -1480 -5770 -1080 -5710
rect -1480 -5850 -1430 -5770
rect -1350 -5850 -1230 -5770
rect -1150 -5850 -1080 -5770
rect -1480 -5870 -1080 -5850
rect 250 -5500 650 -5470
rect 250 -5560 280 -5500
rect 340 -5560 400 -5500
rect 460 -5560 520 -5500
rect 580 -5560 650 -5500
rect 250 -5630 650 -5560
rect 250 -5710 300 -5630
rect 380 -5710 500 -5630
rect 580 -5710 650 -5630
rect 250 -5770 650 -5710
rect 250 -5850 300 -5770
rect 380 -5850 500 -5770
rect 580 -5850 650 -5770
rect 250 -5870 650 -5850
rect 2090 -5500 2490 -5470
rect 2090 -5560 2120 -5500
rect 2180 -5560 2240 -5500
rect 2300 -5560 2360 -5500
rect 2420 -5560 2490 -5500
rect 2090 -5630 2490 -5560
rect 2090 -5710 2140 -5630
rect 2220 -5710 2340 -5630
rect 2420 -5710 2490 -5630
rect 2090 -5770 2490 -5710
rect 9110 -5720 9310 -5110
rect 2090 -5850 2140 -5770
rect 2220 -5850 2340 -5770
rect 2420 -5850 2490 -5770
rect 2090 -5870 2490 -5850
rect 7200 -5920 9310 -5720
rect 7200 -6050 7400 -5920
rect 5020 -6100 7400 -6050
rect 2800 -6110 3200 -6100
rect 2800 -6360 3280 -6110
rect 2800 -6460 2920 -6360
rect 3020 -6460 3120 -6360
rect 3220 -6460 3280 -6360
rect 5020 -6200 5070 -6100
rect 5170 -6200 5270 -6100
rect 5370 -6200 7400 -6100
rect 5020 -6250 7400 -6200
rect 5020 -6310 5220 -6250
rect 5020 -6410 5070 -6310
rect 5170 -6410 5220 -6310
rect 5020 -6460 5220 -6410
rect 2800 -6530 3280 -6460
rect 2800 -6630 3020 -6530
rect 3120 -6630 3280 -6530
rect -1960 -7090 -1480 -7060
rect -1960 -7150 -1930 -7090
rect -1870 -7150 -1810 -7090
rect -1750 -7150 -1690 -7090
rect -1630 -7150 -1570 -7090
rect -1510 -7150 -1480 -7090
rect -1960 -7210 -1480 -7150
rect -1960 -7290 -1930 -7210
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -1960 -7320 -1480 -7290
rect -2800 -7910 -2600 -7860
rect -2800 -7970 -2730 -7910
rect -2670 -7970 -2600 -7910
rect -2800 -8030 -2600 -7970
rect -2800 -8090 -2730 -8030
rect -2670 -8090 -2600 -8030
rect -2800 -8150 -2600 -8090
rect -2800 -8210 -2730 -8150
rect -2670 -8210 -2600 -8150
rect -2800 -8640 -2600 -8210
rect -2800 -8840 -1980 -8640
rect -2380 -24100 -1980 -8840
rect -150 -9160 250 -9140
rect -150 -9220 -120 -9160
rect -60 -9220 0 -9160
rect 60 -9220 120 -9160
rect 180 -9220 250 -9160
rect -150 -9260 250 -9220
rect -150 -9340 -120 -9260
rect -40 -9340 110 -9260
rect 190 -9340 250 -9260
rect -150 -9360 250 -9340
rect -1840 -9570 -1440 -9550
rect -1840 -9630 -1810 -9570
rect -1750 -9630 -1690 -9570
rect -1630 -9630 -1570 -9570
rect -1510 -9630 -1440 -9570
rect -1840 -9660 -1440 -9630
rect -1840 -9740 -1810 -9660
rect -1730 -9740 -1580 -9660
rect -1500 -9740 -1440 -9660
rect -1840 -9770 -1440 -9740
rect -2380 -24500 -790 -24100
rect -1190 -25254 -790 -24500
rect 2800 -25158 3280 -6630
rect 18510 -7010 18760 -6940
rect 18510 -7070 18530 -7010
rect 18590 -7070 18760 -7010
rect 18510 -7130 18650 -7070
rect 18510 -7190 18530 -7130
rect 18590 -7150 18650 -7130
rect 18730 -7150 18760 -7070
rect 18590 -7190 18760 -7150
rect 18510 -7230 18760 -7190
rect 18510 -7250 18650 -7230
rect 18510 -7310 18530 -7250
rect 18590 -7310 18650 -7250
rect 18730 -7310 18760 -7230
rect 18510 -7340 18760 -7310
rect 10000 -9580 10390 -9560
rect 10000 -9640 10030 -9580
rect 10090 -9640 10150 -9580
rect 10210 -9640 10270 -9580
rect 10330 -9640 10390 -9580
rect 10000 -9690 10390 -9640
rect 10000 -9770 10040 -9690
rect 10120 -9770 10260 -9690
rect 10340 -9770 10390 -9690
rect 10000 -9800 10390 -9770
rect 16070 -9580 16460 -9560
rect 16070 -9640 16090 -9580
rect 16150 -9640 16210 -9580
rect 16270 -9640 16330 -9580
rect 16390 -9640 16460 -9580
rect 16070 -9690 16460 -9640
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9800 16460 -9770
rect -7406 -26634 -6946 -25254
rect -1248 -26634 -696 -25254
rect 2800 -26630 3352 -25158
<< via2 >>
rect -670 8100 -590 8180
rect -430 8100 -350 8180
rect 3260 8110 3340 8190
rect 3480 8110 3560 8190
rect 11080 8110 11160 8190
rect 11310 8110 11390 8190
rect 15900 8100 15980 8180
rect 16140 8100 16220 8180
rect 14830 4540 14930 4640
rect 14830 4340 14930 4440
rect -1430 880 -1350 960
rect -1220 880 -1140 960
rect -1430 740 -1350 820
rect -1220 740 -1140 820
rect -270 870 -190 950
rect -50 870 30 950
rect -270 730 -190 810
rect -50 730 30 810
rect 930 900 1010 980
rect 1170 900 1250 980
rect 930 740 1010 820
rect 1170 740 1250 820
rect 4650 -1000 4750 -900
rect 4860 -1000 4960 -900
rect 4860 -1210 4960 -1110
rect 2380 -3420 2460 -3340
rect 2540 -3420 2620 -3340
rect -2290 -4300 -2210 -4220
rect -2040 -4300 -1960 -4220
rect -2290 -4450 -2210 -4370
rect -2040 -4450 -1960 -4370
rect 18650 -2470 18730 -2390
rect 18650 -2630 18730 -2550
rect 13300 -3650 13380 -3570
rect 13300 -3890 13380 -3810
rect -1430 -5710 -1350 -5630
rect -1230 -5710 -1150 -5630
rect -1430 -5850 -1350 -5770
rect -1230 -5850 -1150 -5770
rect 300 -5710 380 -5630
rect 500 -5710 580 -5630
rect 300 -5850 380 -5770
rect 500 -5850 580 -5770
rect 2140 -5710 2220 -5630
rect 2340 -5710 2420 -5630
rect 2140 -5850 2220 -5770
rect 2340 -5850 2420 -5770
rect 5070 -6200 5170 -6100
rect 5270 -6200 5370 -6100
rect 5070 -6410 5170 -6310
rect -1930 -7290 -1850 -7210
rect -1770 -7290 -1690 -7210
rect -1610 -7290 -1530 -7210
rect -120 -9340 -40 -9260
rect 110 -9340 190 -9260
rect -1810 -9740 -1730 -9660
rect -1580 -9740 -1500 -9660
rect 18650 -7150 18730 -7070
rect 18650 -7310 18730 -7230
rect 10040 -9770 10120 -9690
rect 10260 -9770 10340 -9690
rect 16100 -9770 16180 -9690
rect 16340 -9770 16420 -9690
<< metal3 >>
rect -15436 26070 -13804 26452
rect -15436 25670 -10370 26070
rect -15436 25500 -13804 25670
rect -10770 -840 -10370 25670
rect -8930 11810 24960 11960
rect -8930 11740 -670 11810
rect -8930 11640 -8840 11740
rect -8740 11640 -8640 11740
rect -8540 11710 -670 11740
rect -570 11710 -470 11810
rect -370 11780 24960 11810
rect -370 11710 3260 11780
rect -8540 11680 3260 11710
rect 3360 11680 3460 11780
rect 3560 11740 24960 11780
rect 3560 11730 15920 11740
rect 3560 11680 11080 11730
rect -8540 11640 11080 11680
rect -8930 11630 11080 11640
rect 11180 11630 11280 11730
rect 11380 11640 15920 11730
rect 16020 11640 16120 11740
rect 16220 11730 24960 11740
rect 16220 11640 24420 11730
rect 11380 11630 24420 11640
rect 24520 11630 24620 11730
rect 24720 11630 24960 11730
rect -8930 11610 24960 11630
rect -8930 11540 -670 11610
rect -8930 11440 -8840 11540
rect -8740 11440 -8640 11540
rect -8540 11510 -670 11540
rect -570 11510 -470 11610
rect -370 11580 24960 11610
rect -370 11510 3260 11580
rect -8540 11480 3260 11510
rect 3360 11480 3460 11580
rect 3560 11540 24960 11580
rect 3560 11530 15920 11540
rect 3560 11480 11080 11530
rect -8540 11440 11080 11480
rect -8930 11430 11080 11440
rect 11180 11430 11280 11530
rect 11380 11440 15920 11530
rect 16020 11440 16120 11540
rect 16220 11530 24960 11540
rect 16220 11440 24420 11530
rect 11380 11430 24420 11440
rect 24520 11430 24620 11530
rect 24720 11430 24960 11530
rect -8930 11340 24960 11430
rect -4160 9740 20150 9900
rect -4160 9640 -4070 9740
rect -3970 9640 -3870 9740
rect -3770 9730 20150 9740
rect -3770 9640 19700 9730
rect -4160 9630 19700 9640
rect 19800 9630 19900 9730
rect 20000 9630 20150 9730
rect -4160 9540 20150 9630
rect -4160 9440 -4070 9540
rect -3970 9440 -3870 9540
rect -3770 9530 20150 9540
rect -3770 9440 19700 9530
rect -4160 9430 19700 9440
rect 19800 9430 19900 9530
rect 20000 9430 20150 9530
rect -4160 9300 20150 9430
rect -710 8350 -310 8370
rect -710 8250 -670 8350
rect -570 8250 -470 8350
rect -370 8250 -310 8350
rect -710 8200 -310 8250
rect -710 8080 -690 8200
rect -570 8080 -450 8200
rect -330 8080 -310 8200
rect -710 8070 -310 8080
rect 3220 8350 3620 8370
rect 3220 8250 3260 8350
rect 3360 8250 3460 8350
rect 3560 8250 3620 8350
rect 3220 8190 3620 8250
rect 3220 8110 3260 8190
rect 3340 8110 3480 8190
rect 3560 8110 3620 8190
rect 3220 8070 3620 8110
rect 11040 8350 11440 8370
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 8190 11440 8250
rect 11040 8110 11080 8190
rect 11160 8110 11310 8190
rect 11390 8110 11440 8190
rect 11040 8070 11440 8110
rect 15870 8330 16270 8350
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 8180 16270 8230
rect 15870 8100 15900 8180
rect 15980 8100 16140 8180
rect 16220 8100 16270 8180
rect 15870 8070 16270 8100
rect 14680 4640 20150 4700
rect 14680 4540 14830 4640
rect 14930 4540 19700 4640
rect 19800 4540 19900 4640
rect 20000 4540 20150 4640
rect 14680 4440 20150 4540
rect 14680 4340 14830 4440
rect 14930 4340 19700 4440
rect 19800 4340 19900 4440
rect 20000 4340 20150 4440
rect 14680 4300 20150 4340
rect -8930 1050 1290 1110
rect -8930 950 -8850 1050
rect -8750 950 -8650 1050
rect -8550 980 1290 1050
rect -8550 960 930 980
rect -8550 950 -1430 960
rect -8930 880 -1430 950
rect -1350 880 -1220 960
rect -1140 950 930 960
rect -1140 880 -270 950
rect -8930 870 -270 880
rect -190 870 -50 950
rect 30 900 930 950
rect 1010 900 1170 980
rect 1250 900 1290 980
rect 30 870 1290 900
rect -8930 850 1290 870
rect -8930 750 -8850 850
rect -8750 750 -8650 850
rect -8550 820 1290 850
rect -8550 750 -1430 820
rect -8930 740 -1430 750
rect -1350 740 -1220 820
rect -1140 810 930 820
rect -1140 740 -270 810
rect -8930 730 -270 740
rect -190 730 -50 810
rect 30 740 930 810
rect 1010 740 1170 820
rect 1250 740 1290 820
rect 30 730 1290 740
rect -8930 710 1290 730
rect -10770 -900 5020 -840
rect -10770 -1000 4650 -900
rect 4750 -1000 4860 -900
rect 4960 -1000 5020 -900
rect -10770 -1060 5020 -1000
rect 4800 -1110 5020 -1060
rect 4800 -1210 4860 -1110
rect 4960 -1210 5020 -1110
rect 4800 -1250 5020 -1210
rect 18510 -2390 20150 -2340
rect 18510 -2470 18650 -2390
rect 18730 -2470 19710 -2390
rect 18510 -2490 19710 -2470
rect 19810 -2490 19910 -2390
rect 20010 -2490 20150 -2390
rect 18510 -2550 20150 -2490
rect 18510 -2630 18650 -2550
rect 18730 -2590 20150 -2550
rect 18730 -2630 19710 -2590
rect 18510 -2690 19710 -2630
rect 19810 -2690 19910 -2590
rect 20010 -2690 20150 -2590
rect 18510 -2740 20150 -2690
rect -4130 -3120 2760 -3080
rect -4130 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 2760 -3120
rect -4130 -3320 2760 -3220
rect -4130 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3340 2760 -3320
rect -3770 -3420 2380 -3340
rect 2460 -3420 2540 -3340
rect 2620 -3420 2760 -3340
rect -4130 -3480 2760 -3420
rect 13160 -3570 24960 -3540
rect 13160 -3650 13300 -3570
rect 13380 -3580 24960 -3570
rect 13380 -3650 24430 -3580
rect 13160 -3680 24430 -3650
rect 24530 -3680 24630 -3580
rect 24730 -3680 24960 -3580
rect 13160 -3780 24960 -3680
rect 13160 -3810 24430 -3780
rect 13160 -3890 13300 -3810
rect 13380 -3880 24430 -3810
rect 24530 -3880 24630 -3780
rect 24730 -3880 24960 -3780
rect 13380 -3890 24960 -3880
rect 13160 -3930 24960 -3890
rect 13160 -3940 23950 -3930
rect -8930 -4220 -1920 -4190
rect -8930 -4230 -2290 -4220
rect -8930 -4330 -8840 -4230
rect -8740 -4330 -8640 -4230
rect -8540 -4300 -2290 -4230
rect -2210 -4300 -2040 -4220
rect -1960 -4300 -1920 -4220
rect -8540 -4330 -1920 -4300
rect -8930 -4370 -1920 -4330
rect -8930 -4430 -2290 -4370
rect -8930 -4530 -8840 -4430
rect -8740 -4530 -8640 -4430
rect -8540 -4450 -2290 -4430
rect -2210 -4450 -2040 -4370
rect -1960 -4450 -1920 -4370
rect -8540 -4530 -1920 -4450
rect -8930 -4590 -1920 -4530
rect -3290 -5630 2490 -5470
rect -3290 -5710 -1430 -5630
rect -1350 -5710 -1230 -5630
rect -1150 -5710 300 -5630
rect 380 -5710 500 -5630
rect 580 -5710 2140 -5630
rect 2220 -5710 2340 -5630
rect 2420 -5710 2490 -5630
rect -3290 -5770 2490 -5710
rect -3290 -5850 -1430 -5770
rect -1350 -5850 -1230 -5770
rect -1150 -5850 300 -5770
rect 380 -5850 500 -5770
rect 580 -5850 2140 -5770
rect 2220 -5850 2340 -5770
rect 2420 -5850 2490 -5770
rect -3290 -5870 2490 -5850
rect -3290 -6260 -2870 -5870
rect 5220 -6050 5420 -6040
rect -3450 -6270 -2870 -6260
rect -4130 -6320 -2870 -6270
rect -4130 -6420 -4090 -6320
rect -3990 -6420 -3890 -6320
rect -3790 -6420 -2870 -6320
rect -4130 -6520 -2870 -6420
rect -4130 -6620 -4090 -6520
rect -3990 -6620 -3890 -6520
rect -3790 -6620 -2870 -6520
rect -4130 -6670 -2870 -6620
rect 5020 -6100 5420 -6050
rect 5020 -6200 5070 -6100
rect 5170 -6200 5270 -6100
rect 5370 -6200 5420 -6100
rect 5020 -6250 5420 -6200
rect 5020 -6310 5220 -6250
rect 5020 -6410 5070 -6310
rect 5170 -6410 5220 -6310
rect -4130 -7080 -1480 -7030
rect -4130 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -1480 -7080
rect -4130 -7210 -1480 -7180
rect -4130 -7280 -1930 -7210
rect -4130 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7290 -1930 -7280
rect -1850 -7290 -1770 -7210
rect -1690 -7290 -1610 -7210
rect -1530 -7290 -1480 -7210
rect -3790 -7320 -1480 -7290
rect -3790 -7380 -3600 -7320
rect -4130 -7430 -3600 -7380
rect -150 -9260 250 -9240
rect -150 -9340 -120 -9260
rect -40 -9340 110 -9260
rect 190 -9340 250 -9260
rect -150 -9370 250 -9340
rect -150 -9470 -130 -9370
rect -30 -9470 70 -9370
rect 170 -9470 250 -9370
rect -150 -9480 250 -9470
rect -1840 -9660 -1440 -9640
rect -1840 -9740 -1810 -9660
rect -1730 -9740 -1580 -9660
rect -1500 -9740 -1440 -9660
rect -1840 -9780 -1440 -9740
rect -1840 -9880 -1810 -9780
rect -1710 -9880 -1610 -9780
rect -1510 -9880 -1440 -9780
rect -1840 -9900 -1440 -9880
rect 5020 -11700 5220 -6410
rect 18510 -6990 20150 -6940
rect 18510 -7070 19700 -6990
rect 18510 -7150 18650 -7070
rect 18730 -7090 19700 -7070
rect 19800 -7090 19900 -6990
rect 20000 -7090 20150 -6990
rect 18730 -7150 20150 -7090
rect 18510 -7190 20150 -7150
rect 18510 -7230 19700 -7190
rect 18510 -7310 18650 -7230
rect 18730 -7290 19700 -7230
rect 19800 -7290 19900 -7190
rect 20000 -7290 20150 -7190
rect 18730 -7310 20150 -7290
rect 18510 -7340 20150 -7310
rect 10000 -9690 10390 -9660
rect 10000 -9770 10040 -9690
rect 10120 -9770 10260 -9690
rect 10340 -9770 10390 -9690
rect 10000 -9800 10390 -9770
rect 10000 -9900 10030 -9800
rect 10130 -9900 10250 -9800
rect 10350 -9900 10390 -9800
rect 10000 -9910 10390 -9900
rect 16070 -9690 16460 -9660
rect 16070 -9770 16100 -9690
rect 16180 -9770 16340 -9690
rect 16420 -9770 16460 -9690
rect 16070 -9820 16460 -9770
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -9940 16460 -9920
rect -12420 -11900 5220 -11700
rect -15436 -26170 -13804 -25772
rect -12420 -26170 -12020 -11900
rect -4160 -18710 20150 -18500
rect -4160 -18810 -4070 -18710
rect -3970 -18810 -3870 -18710
rect -3770 -18720 20150 -18710
rect -3770 -18810 10040 -18720
rect -4160 -18820 10040 -18810
rect 10140 -18820 10240 -18720
rect 10340 -18820 16120 -18720
rect 16220 -18820 16320 -18720
rect 16420 -18730 20150 -18720
rect 16420 -18820 19690 -18730
rect -4160 -18830 19690 -18820
rect 19790 -18830 19890 -18730
rect 19990 -18830 20150 -18730
rect -4160 -18910 20150 -18830
rect -4160 -19010 -4070 -18910
rect -3970 -19010 -3870 -18910
rect -3770 -18920 20150 -18910
rect -3770 -19010 10040 -18920
rect -4160 -19020 10040 -19010
rect 10140 -19020 10240 -18920
rect 10340 -19020 16120 -18920
rect 16220 -19020 16320 -18920
rect 16420 -18930 20150 -18920
rect 16420 -19020 19690 -18930
rect -4160 -19030 19690 -19020
rect 19790 -19030 19890 -18930
rect 19990 -19030 20150 -18930
rect -4160 -19120 20150 -19030
rect -8930 -23090 24960 -22880
rect -8930 -23120 -1800 -23090
rect -8930 -23220 -8840 -23120
rect -8740 -23220 -8640 -23120
rect -8540 -23190 -1800 -23120
rect -1700 -23190 -1600 -23090
rect -1500 -23110 24960 -23090
rect -1500 -23190 -100 -23110
rect -8540 -23210 -100 -23190
rect 0 -23210 100 -23110
rect 200 -23130 24960 -23110
rect 200 -23210 24420 -23130
rect -8540 -23220 24420 -23210
rect -8930 -23230 24420 -23220
rect 24520 -23230 24620 -23130
rect 24720 -23230 24960 -23130
rect -8930 -23290 24960 -23230
rect -8930 -23320 -1800 -23290
rect -8930 -23420 -8840 -23320
rect -8740 -23420 -8640 -23320
rect -8540 -23390 -1800 -23320
rect -1700 -23390 -1600 -23290
rect -1500 -23310 24960 -23290
rect -1500 -23390 -100 -23310
rect -8540 -23410 -100 -23390
rect 0 -23410 100 -23310
rect 200 -23330 24960 -23310
rect 200 -23410 24420 -23330
rect -8540 -23420 24420 -23410
rect -8930 -23430 24420 -23420
rect 24520 -23430 24620 -23330
rect 24720 -23430 24960 -23330
rect -8930 -23480 24960 -23430
rect -15436 -26570 -12020 -26170
rect -15436 -26724 -13804 -26570
<< via3 >>
rect -8840 11640 -8740 11740
rect -8640 11640 -8540 11740
rect -670 11710 -570 11810
rect -470 11710 -370 11810
rect 3260 11680 3360 11780
rect 3460 11680 3560 11780
rect 11080 11630 11180 11730
rect 11280 11630 11380 11730
rect 15920 11640 16020 11740
rect 16120 11640 16220 11740
rect 24420 11630 24520 11730
rect 24620 11630 24720 11730
rect -8840 11440 -8740 11540
rect -8640 11440 -8540 11540
rect -670 11510 -570 11610
rect -470 11510 -370 11610
rect 3260 11480 3360 11580
rect 3460 11480 3560 11580
rect 11080 11430 11180 11530
rect 11280 11430 11380 11530
rect 15920 11440 16020 11540
rect 16120 11440 16220 11540
rect 24420 11430 24520 11530
rect 24620 11430 24720 11530
rect -4070 9640 -3970 9740
rect -3870 9640 -3770 9740
rect 19700 9630 19800 9730
rect 19900 9630 20000 9730
rect -4070 9440 -3970 9540
rect -3870 9440 -3770 9540
rect 19700 9430 19800 9530
rect 19900 9430 20000 9530
rect -670 8250 -570 8350
rect -470 8250 -370 8350
rect -690 8180 -570 8200
rect -690 8100 -670 8180
rect -670 8100 -590 8180
rect -590 8100 -570 8180
rect -690 8080 -570 8100
rect -450 8180 -330 8200
rect -450 8100 -430 8180
rect -430 8100 -350 8180
rect -350 8100 -330 8180
rect -450 8080 -330 8100
rect 3260 8250 3360 8350
rect 3460 8250 3560 8350
rect 11080 8250 11180 8350
rect 11280 8250 11380 8350
rect 15900 8230 16000 8330
rect 16130 8230 16230 8330
rect 19700 4540 19800 4640
rect 19900 4540 20000 4640
rect 19700 4340 19800 4440
rect 19900 4340 20000 4440
rect -8850 950 -8750 1050
rect -8650 950 -8550 1050
rect -8850 750 -8750 850
rect -8650 750 -8550 850
rect 19710 -2490 19810 -2390
rect 19910 -2490 20010 -2390
rect 19710 -2690 19810 -2590
rect 19910 -2690 20010 -2590
rect -4070 -3220 -3970 -3120
rect -3870 -3220 -3770 -3120
rect -4070 -3420 -3970 -3320
rect -3870 -3420 -3770 -3320
rect 24430 -3680 24530 -3580
rect 24630 -3680 24730 -3580
rect 24430 -3880 24530 -3780
rect 24630 -3880 24730 -3780
rect -8840 -4330 -8740 -4230
rect -8640 -4330 -8540 -4230
rect -8840 -4530 -8740 -4430
rect -8640 -4530 -8540 -4430
rect -4090 -6420 -3990 -6320
rect -3890 -6420 -3790 -6320
rect -4090 -6620 -3990 -6520
rect -3890 -6620 -3790 -6520
rect -4090 -7180 -3990 -7080
rect -3890 -7180 -3790 -7080
rect -4090 -7380 -3990 -7280
rect -3890 -7380 -3790 -7280
rect -130 -9470 -30 -9370
rect 70 -9470 170 -9370
rect -1810 -9880 -1710 -9780
rect -1610 -9880 -1510 -9780
rect 19700 -7090 19800 -6990
rect 19900 -7090 20000 -6990
rect 19700 -7290 19800 -7190
rect 19900 -7290 20000 -7190
rect 10030 -9900 10130 -9800
rect 10250 -9900 10350 -9800
rect 16110 -9920 16210 -9820
rect 16310 -9920 16410 -9820
rect -4070 -18810 -3970 -18710
rect -3870 -18810 -3770 -18710
rect 10040 -18820 10140 -18720
rect 10240 -18820 10340 -18720
rect 16120 -18820 16220 -18720
rect 16320 -18820 16420 -18720
rect 19690 -18830 19790 -18730
rect 19890 -18830 19990 -18730
rect -4070 -19010 -3970 -18910
rect -3870 -19010 -3770 -18910
rect 10040 -19020 10140 -18920
rect 10240 -19020 10340 -18920
rect 16120 -19020 16220 -18920
rect 16320 -19020 16420 -18920
rect 19690 -19030 19790 -18930
rect 19890 -19030 19990 -18930
rect -8840 -23220 -8740 -23120
rect -8640 -23220 -8540 -23120
rect -1800 -23190 -1700 -23090
rect -1600 -23190 -1500 -23090
rect -100 -23210 0 -23110
rect 100 -23210 200 -23110
rect 24420 -23230 24520 -23130
rect 24620 -23230 24720 -23130
rect -8840 -23420 -8740 -23320
rect -8640 -23420 -8540 -23320
rect -1800 -23390 -1700 -23290
rect -1600 -23390 -1500 -23290
rect -100 -23410 0 -23310
rect 100 -23410 200 -23310
rect 24420 -23430 24520 -23330
rect 24620 -23430 24720 -23330
<< metal4 >>
rect -8930 11740 -8310 11960
rect -8930 11640 -8840 11740
rect -8740 11640 -8640 11740
rect -8540 11640 -8310 11740
rect -8930 11540 -8310 11640
rect -8930 11440 -8840 11540
rect -8740 11440 -8640 11540
rect -8540 11440 -8310 11540
rect -8930 1050 -8310 11440
rect -710 11810 -310 11960
rect -710 11710 -670 11810
rect -570 11710 -470 11810
rect -370 11710 -310 11810
rect -710 11610 -310 11710
rect -710 11510 -670 11610
rect -570 11510 -470 11610
rect -370 11510 -310 11610
rect -8930 950 -8850 1050
rect -8750 950 -8650 1050
rect -8550 950 -8310 1050
rect -8930 850 -8310 950
rect -8930 750 -8850 850
rect -8750 750 -8650 850
rect -8550 750 -8310 850
rect -8930 -4230 -8310 750
rect -8930 -4330 -8840 -4230
rect -8740 -4330 -8640 -4230
rect -8540 -4330 -8310 -4230
rect -8930 -4430 -8310 -4330
rect -8930 -4530 -8840 -4430
rect -8740 -4530 -8640 -4430
rect -8540 -4530 -8310 -4430
rect -8930 -23120 -8310 -4530
rect -4160 9740 -3560 9900
rect -4160 9640 -4070 9740
rect -3970 9640 -3870 9740
rect -3770 9640 -3560 9740
rect -4160 9540 -3560 9640
rect -4160 9440 -4070 9540
rect -3970 9440 -3870 9540
rect -3770 9440 -3560 9540
rect -4160 -3120 -3560 9440
rect -710 8350 -310 11510
rect -710 8250 -670 8350
rect -570 8250 -470 8350
rect -370 8250 -310 8350
rect -710 8200 -310 8250
rect -710 8080 -690 8200
rect -570 8080 -450 8200
rect -330 8080 -310 8200
rect -710 7990 -310 8080
rect 3220 11780 3620 11960
rect 3220 11680 3260 11780
rect 3360 11680 3460 11780
rect 3560 11680 3620 11780
rect 3220 11580 3620 11680
rect 3220 11480 3260 11580
rect 3360 11480 3460 11580
rect 3560 11480 3620 11580
rect 3220 8350 3620 11480
rect 3220 8250 3260 8350
rect 3360 8250 3460 8350
rect 3560 8250 3620 8350
rect 3220 7990 3620 8250
rect 11040 11730 11440 11960
rect 11040 11630 11080 11730
rect 11180 11630 11280 11730
rect 11380 11630 11440 11730
rect 11040 11530 11440 11630
rect 11040 11430 11080 11530
rect 11180 11430 11280 11530
rect 11380 11430 11440 11530
rect 11040 8350 11440 11430
rect 11040 8250 11080 8350
rect 11180 8250 11280 8350
rect 11380 8250 11440 8350
rect 11040 7990 11440 8250
rect 15870 11740 16270 11960
rect 24360 11900 24960 11960
rect 15870 11640 15920 11740
rect 16020 11640 16120 11740
rect 16220 11640 16270 11740
rect 15870 11540 16270 11640
rect 15870 11440 15920 11540
rect 16020 11440 16120 11540
rect 16220 11440 16270 11540
rect 15870 8330 16270 11440
rect 24356 11730 24960 11900
rect 24356 11630 24420 11730
rect 24520 11630 24620 11730
rect 24720 11630 24960 11730
rect 24356 11530 24960 11630
rect 24356 11430 24420 11530
rect 24520 11430 24620 11530
rect 24720 11430 24960 11530
rect 19520 9860 20150 9900
rect 15870 8230 15900 8330
rect 16000 8230 16130 8330
rect 16230 8230 16270 8330
rect 15870 7990 16270 8230
rect 19516 9730 20150 9860
rect 19516 9630 19700 9730
rect 19800 9630 19900 9730
rect 20000 9630 20150 9730
rect 19516 9530 20150 9630
rect 19516 9430 19700 9530
rect 19800 9430 19900 9530
rect 20000 9430 20150 9530
rect -4160 -3220 -4070 -3120
rect -3970 -3220 -3870 -3120
rect -3770 -3220 -3560 -3120
rect -4160 -3320 -3560 -3220
rect -4160 -3420 -4070 -3320
rect -3970 -3420 -3870 -3320
rect -3770 -3420 -3560 -3320
rect -4160 -6320 -3560 -3420
rect -4160 -6420 -4090 -6320
rect -3990 -6420 -3890 -6320
rect -3790 -6420 -3560 -6320
rect -4160 -6520 -3560 -6420
rect -4160 -6620 -4090 -6520
rect -3990 -6620 -3890 -6520
rect -3790 -6620 -3560 -6520
rect -4160 -7080 -3560 -6620
rect -4160 -7180 -4090 -7080
rect -3990 -7180 -3890 -7080
rect -3790 -7180 -3560 -7080
rect -4160 -7280 -3560 -7180
rect -4160 -7380 -4090 -7280
rect -3990 -7380 -3890 -7280
rect -3790 -7380 -3560 -7280
rect -4160 -18710 -3560 -7380
rect 19516 4640 20150 9430
rect 19516 4540 19700 4640
rect 19800 4540 19900 4640
rect 20000 4540 20150 4640
rect 19516 4440 20150 4540
rect 19516 4340 19700 4440
rect 19800 4340 19900 4440
rect 20000 4340 20150 4440
rect 19516 -2390 20150 4340
rect 19516 -2490 19710 -2390
rect 19810 -2490 19910 -2390
rect 20010 -2490 20150 -2390
rect 19516 -2590 20150 -2490
rect 19516 -2690 19710 -2590
rect 19810 -2690 19910 -2590
rect 20010 -2690 20150 -2590
rect 19516 -6990 20150 -2690
rect 19516 -7090 19700 -6990
rect 19800 -7090 19900 -6990
rect 20000 -7090 20150 -6990
rect 19516 -7190 20150 -7090
rect 19516 -7290 19700 -7190
rect 19800 -7290 19900 -7190
rect 20000 -7290 20150 -7190
rect -150 -9370 250 -9140
rect -150 -9470 -130 -9370
rect -30 -9470 70 -9370
rect 170 -9470 250 -9370
rect -4160 -18810 -4070 -18710
rect -3970 -18810 -3870 -18710
rect -3770 -18810 -3560 -18710
rect -4160 -18910 -3560 -18810
rect -4160 -19010 -4070 -18910
rect -3970 -19010 -3870 -18910
rect -3770 -19010 -3560 -18910
rect -4160 -19120 -3560 -19010
rect -1840 -9780 -1440 -9550
rect -1840 -9880 -1810 -9780
rect -1710 -9880 -1610 -9780
rect -1510 -9880 -1440 -9780
rect -8930 -23220 -8840 -23120
rect -8740 -23220 -8640 -23120
rect -8540 -23220 -8310 -23120
rect -8930 -23320 -8310 -23220
rect -8930 -23420 -8840 -23320
rect -8740 -23420 -8640 -23320
rect -8540 -23420 -8310 -23320
rect -8930 -23480 -8310 -23420
rect -1840 -23090 -1440 -9880
rect -1840 -23190 -1800 -23090
rect -1700 -23190 -1600 -23090
rect -1500 -23190 -1440 -23090
rect -1840 -23290 -1440 -23190
rect -1840 -23390 -1800 -23290
rect -1700 -23390 -1600 -23290
rect -1500 -23390 -1440 -23290
rect -1840 -23480 -1440 -23390
rect -150 -23110 250 -9470
rect 10000 -9800 10390 -9550
rect 10000 -9900 10030 -9800
rect 10130 -9900 10250 -9800
rect 10350 -9900 10390 -9800
rect 10000 -18720 10390 -9900
rect 10000 -18820 10040 -18720
rect 10140 -18820 10240 -18720
rect 10340 -18820 10390 -18720
rect 10000 -18920 10390 -18820
rect 10000 -19020 10040 -18920
rect 10140 -19020 10240 -18920
rect 10340 -19020 10390 -18920
rect 10000 -19115 10390 -19020
rect 16070 -9820 16460 -9560
rect 16070 -9920 16110 -9820
rect 16210 -9920 16310 -9820
rect 16410 -9920 16460 -9820
rect 16070 -18720 16460 -9920
rect 16070 -18820 16120 -18720
rect 16220 -18820 16320 -18720
rect 16420 -18820 16460 -18720
rect 16070 -18920 16460 -18820
rect 16070 -19020 16120 -18920
rect 16220 -19020 16320 -18920
rect 16420 -19020 16460 -18920
rect 16070 -19115 16460 -19020
rect 19516 -18730 20150 -7290
rect 19516 -18830 19690 -18730
rect 19790 -18830 19890 -18730
rect 19990 -18830 20150 -18730
rect 19516 -18930 20150 -18830
rect 19516 -19030 19690 -18930
rect 19790 -19030 19890 -18930
rect 19990 -19030 20150 -18930
rect 19516 -19100 20150 -19030
rect 19520 -19120 20150 -19100
rect 24356 -3580 24960 11430
rect 24356 -3680 24430 -3580
rect 24530 -3680 24630 -3580
rect 24730 -3680 24960 -3580
rect 24356 -3780 24960 -3680
rect 24356 -3880 24430 -3780
rect 24530 -3880 24630 -3780
rect 24730 -3880 24960 -3780
rect -150 -23210 -100 -23110
rect 0 -23210 100 -23110
rect 200 -23210 250 -23110
rect -150 -23310 250 -23210
rect -150 -23410 -100 -23310
rect 0 -23410 100 -23310
rect 200 -23410 250 -23310
rect -150 -23470 250 -23410
rect 24356 -23130 24960 -3880
rect 24356 -23230 24420 -23130
rect 24520 -23230 24620 -23130
rect 24720 -23230 24960 -23130
rect 24356 -23330 24960 -23230
rect 24356 -23430 24420 -23330
rect 24520 -23430 24620 -23330
rect 24720 -23430 24960 -23330
rect 24356 -23476 24960 -23430
rect 24360 -23480 24960 -23476
use ALib_DCO  ALib_DCO_0
timestamp 1731453370
transform 1 0 5200 0 1 -5190
box 1000 -4470 13410 5980
use ALib_VCO  ALib_VCO_0
timestamp 1731453370
transform 1 0 -2020 0 1 1040
box 0 280 20640 7030
use DLib_Quantizer  DLib_Quantizer_0
timestamp 1731453370
transform 1 0 -2210 0 1 -4630
box 190 -710 5890 730
use DLib_UpDownCounter  DLib_UpDownCounter_0
timestamp 1731453370
transform 1 0 -1140 0 1 -5986
box -880 -3154 3140 -440
use DLib_UpDownCounter  DLib_UpDownCounter_1
timestamp 1731453370
transform 1 0 -1140 0 1 344
box -880 -3154 3140 -440
<< labels >>
flabel metal3 -15436 25500 -13804 26452 1 FreeSans 1088 0 0 0 vbias_12
port 1 nsew signal input
flabel metal3 -15436 -26724 -13804 -25772 1 FreeSans 1088 0 0 0 vbias_34
port 2 nsew signal input
flabel metal2 -7406 -26634 -6946 -25254 1 FreeSans 736 0 0 0 clk
port 5 nsew signal input
flabel metal2 2800 -26630 3352 -25158 1 FreeSans 736 0 0 0 quantizer_out
port 6 nsew signal output
flabel metal2 -1248 -26634 -696 -25254 1 FreeSans 736 0 0 0 enable_in
port 4 nsew signal input
flabel metal2 39514 32062 41630 32430 1 FreeSans 1472 0 0 0 analog_in
port 3 nsew signal input
flabel metal4 -8908 -23460 -8364 11900 1 FreeSans 4352 0 0 0 vdda1
port 7 nsew power bidirectional
flabel metal4 -4148 -19108 -3604 9860 1 FreeSans 4352 0 0 0 vssa1
port 8 nsew ground bidirectional
flabel metal3 -4148 -19108 20060 -18564 1 FreeSans 4352 0 0 0 vssa1
port 8 nsew ground bidirectional
flabel metal3 -8908 -23460 24956 -22916 1 FreeSans 4352 0 0 0 vdda1
port 7 nsew power bidirectional
flabel metal3 -8908 11356 24956 11900 1 FreeSans 4352 0 0 0 vdda1
port 7 nsew power bidirectional
flabel metal3 -4148 9316 20060 9860 1 FreeSans 4352 0 0 0 vssa1
port 8 nsew ground bidirectional
<< end >>
