magic
tech sky130A
magscale 1 2
timestamp 1731061822
<< nwell >>
rect 1066 116677 118902 117243
rect 1066 115589 118902 116155
rect 1066 114501 118902 115067
rect 1066 113413 118902 113979
rect 1066 112325 118902 112891
rect 1066 111237 118902 111803
rect 1066 110149 118902 110715
rect 1066 109061 118902 109627
rect 1066 107973 118902 108539
rect 1066 106885 118902 107451
rect 1066 105797 118902 106363
rect 1066 104709 118902 105275
rect 1066 103621 118902 104187
rect 1066 102533 118902 103099
rect 1066 101445 118902 102011
rect 1066 100357 118902 100923
rect 1066 99269 118902 99835
rect 1066 98181 118902 98747
rect 1066 97093 118902 97659
rect 1066 96005 118902 96571
rect 1066 94917 118902 95483
rect 1066 93829 118902 94395
rect 1066 92741 118902 93307
rect 1066 91653 118902 92219
rect 1066 90565 118902 91131
rect 1066 89477 118902 90043
rect 1066 88389 118902 88955
rect 1066 87301 118902 87867
rect 1066 86213 118902 86779
rect 1066 85125 118902 85691
rect 1066 84037 118902 84603
rect 1066 82949 118902 83515
rect 1066 81861 118902 82427
rect 1066 80773 118902 81339
rect 1066 79685 118902 80251
rect 1066 78597 118902 79163
rect 1066 77509 118902 78075
rect 1066 76421 118902 76987
rect 1066 75333 118902 75899
rect 1066 74245 118902 74811
rect 1066 73157 118902 73723
rect 1066 72069 118902 72635
rect 1066 70981 118902 71547
rect 1066 69893 118902 70459
rect 1066 68805 118902 69371
rect 1066 67717 118902 68283
rect 1066 66629 118902 67195
rect 1066 65541 118902 66107
rect 1066 64453 118902 65019
rect 1066 63365 118902 63931
rect 1066 62277 118902 62843
rect 1066 61189 118902 61755
rect 1066 60101 118902 60667
rect 1066 59013 118902 59579
rect 1066 57925 118902 58491
rect 1066 56837 118902 57403
rect 1066 55749 118902 56315
rect 1066 54661 118902 55227
rect 1066 53573 118902 54139
rect 1066 52485 118902 53051
rect 1066 51397 118902 51963
rect 1066 50309 118902 50875
rect 1066 49221 118902 49787
rect 1066 48133 118902 48699
rect 1066 47045 118902 47611
rect 1066 45957 118902 46523
rect 1066 44869 118902 45435
rect 1066 43781 118902 44347
rect 1066 42693 118902 43259
rect 1066 41605 118902 42171
rect 1066 40517 118902 41083
rect 1066 39429 118902 39995
rect 1066 38341 118902 38907
rect 1066 37253 118902 37819
rect 1066 36165 118902 36731
rect 1066 35077 118902 35643
rect 1066 33989 118902 34555
rect 1066 32901 118902 33467
rect 1066 31813 118902 32379
rect 1066 30725 118902 31291
rect 1066 29637 118902 30203
rect 1066 28549 118902 29115
rect 1066 27461 118902 28027
rect 1066 26373 118902 26939
rect 1066 25285 118902 25851
rect 1066 24197 118902 24763
rect 1066 23109 118902 23675
rect 1066 22021 118902 22587
rect 1066 20933 118902 21499
rect 1066 19845 118902 20411
rect 1066 18757 118902 19323
rect 1066 17669 118902 18235
rect 1066 16581 118902 17147
rect 1066 15493 118902 16059
rect 1066 14405 118902 14971
rect 1066 13317 118902 13883
rect 1066 12229 118902 12795
rect 1066 11141 118902 11707
rect 1066 10053 118902 10619
rect 1066 8965 118902 9531
rect 1066 7877 118902 8443
rect 1066 6789 118902 7355
rect 1066 5701 118902 6267
rect 1066 4613 118902 5179
rect 1066 3525 118902 4091
rect 1066 2437 118902 3003
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 1104 2128 118924 117552
<< metal2 >>
rect 6090 119200 6146 120000
rect 18050 119200 18106 120000
rect 30010 119200 30066 120000
rect 41970 119200 42026 120000
rect 53930 119200 53986 120000
rect 65890 119200 65946 120000
rect 77850 119200 77906 120000
rect 89810 119200 89866 120000
rect 101770 119200 101826 120000
rect 113730 119200 113786 120000
<< obsm2 >>
rect 1400 119144 6034 119354
rect 6202 119144 17994 119354
rect 18162 119144 29954 119354
rect 30122 119144 41914 119354
rect 42082 119144 53874 119354
rect 54042 119144 65834 119354
rect 66002 119144 77794 119354
rect 77962 119144 89754 119354
rect 89922 119144 101714 119354
rect 101882 119144 113674 119354
rect 113842 119144 118846 119354
rect 1400 2139 118846 119144
<< metal3 >>
rect 119200 113704 120000 113824
rect 119200 103912 120000 104032
rect 119200 94120 120000 94240
rect 119200 84328 120000 84448
rect 119200 74536 120000 74656
rect 119200 64744 120000 64864
rect 119200 54952 120000 55072
rect 119200 45160 120000 45280
rect 119200 35368 120000 35488
rect 119200 25576 120000 25696
rect 119200 15784 120000 15904
rect 119200 5992 120000 6112
<< obsm3 >>
rect 2129 113904 119200 117537
rect 2129 113624 119120 113904
rect 2129 104112 119200 113624
rect 2129 103832 119120 104112
rect 2129 94320 119200 103832
rect 2129 94040 119120 94320
rect 2129 84528 119200 94040
rect 2129 84248 119120 84528
rect 2129 74736 119200 84248
rect 2129 74456 119120 74736
rect 2129 64944 119200 74456
rect 2129 64664 119120 64944
rect 2129 55152 119200 64664
rect 2129 54872 119120 55152
rect 2129 45360 119200 54872
rect 2129 45080 119120 45360
rect 2129 35568 119200 45080
rect 2129 35288 119120 35568
rect 2129 25776 119200 35288
rect 2129 25496 119120 25776
rect 2129 15984 119200 25496
rect 2129 15704 119120 15984
rect 2129 6192 119200 15704
rect 2129 5912 119120 6192
rect 2129 2143 119200 5912
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 2267 5475 4128 114613
rect 4608 5475 19488 114613
rect 19968 5475 34848 114613
rect 35328 5475 50208 114613
rect 50688 5475 65568 114613
rect 66048 5475 80928 114613
rect 81408 5475 96288 114613
rect 96768 5475 111648 114613
rect 112128 5475 115125 114613
<< labels >>
rlabel metal2 s 89810 119200 89866 120000 6 clk
port 1 nsew signal input
rlabel metal3 s 119200 113704 120000 113824 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 119200 94120 120000 94240 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 119200 74536 120000 74656 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 119200 54952 120000 55072 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 119200 35368 120000 35488 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 119200 15784 120000 15904 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[0]
port 8 nsew signal output
rlabel metal2 s 77850 119200 77906 120000 6 io_oeb[10]
port 9 nsew signal output
rlabel metal2 s 30010 119200 30066 120000 6 io_oeb[1]
port 10 nsew signal output
rlabel metal2 s 6090 119200 6146 120000 6 io_oeb[2]
port 11 nsew signal output
rlabel metal3 s 119200 103912 120000 104032 6 io_oeb[3]
port 12 nsew signal output
rlabel metal3 s 119200 84328 120000 84448 6 io_oeb[4]
port 13 nsew signal output
rlabel metal3 s 119200 64744 120000 64864 6 io_oeb[5]
port 14 nsew signal output
rlabel metal3 s 119200 45160 120000 45280 6 io_oeb[6]
port 15 nsew signal output
rlabel metal3 s 119200 25576 120000 25696 6 io_oeb[7]
port 16 nsew signal output
rlabel metal3 s 119200 5992 120000 6112 6 io_oeb[8]
port 17 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 io_oeb[9]
port 18 nsew signal output
rlabel metal2 s 65890 119200 65946 120000 6 io_out[0]
port 19 nsew signal output
rlabel metal2 s 41970 119200 42026 120000 6 io_out[1]
port 20 nsew signal output
rlabel metal2 s 18050 119200 18106 120000 6 io_out[2]
port 21 nsew signal output
rlabel metal2 s 113730 119200 113786 120000 6 rst
port 22 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 24 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44778336
string GDS_FILE /home/admin/projects/IC5-CASS-2024_2/openlane/hs_ascon/runs/24_11_08_16_06/results/signoff/ascon_wrapper.magic.gds
string GDS_START 901448
<< end >>

