magic
tech sky130A
timestamp 1731473513
<< locali >>
rect 1459 920 1604 960
rect 3036 920 3197 960
rect 4540 950 4580 960
rect 4540 925 4550 950
rect 4575 925 4580 950
rect 4540 920 4580 925
rect 1500 120 1635 130
rect 1465 90 1635 120
rect 3060 90 3215 130
rect 1465 -330 1505 90
rect 2920 -310 3145 -270
rect 4505 -330 4545 110
rect 2922 -1140 3058 -1100
rect 4505 -1105 4545 -1100
rect 4530 -1130 4545 -1105
rect 4505 -1140 4545 -1130
<< viali >>
rect 4550 925 4575 950
rect 4625 925 4650 950
rect 4440 -1130 4465 -1105
rect 4505 -1130 4530 -1105
<< metal1 >>
rect 4540 950 5240 960
rect 4540 925 4550 950
rect 4575 925 4625 950
rect 4650 925 5240 950
rect 4540 920 5240 925
rect -250 670 0 710
rect 4680 670 5090 710
rect -250 -850 -200 670
rect -100 300 0 340
rect 4675 300 4940 340
rect -100 -480 -50 300
rect 4890 -480 4940 300
rect -100 -520 1445 -480
rect 4560 -520 4940 -480
rect 5040 -850 5090 670
rect -250 -890 1445 -850
rect 4530 -890 5090 -850
rect 5190 -1100 5240 920
rect 4425 -1105 5240 -1100
rect 4425 -1130 4440 -1105
rect 4465 -1130 4505 -1105
rect 4530 -1130 5240 -1105
rect 4425 -1140 5240 -1130
use cc_inv_dco  cc_inv_dco_0
timestamp 1730452893
transform 1 0 0 0 1 90
box 0 0 1560 870
use cc_inv_dco  cc_inv_dco_1
timestamp 1730452893
transform 1 0 1560 0 1 90
box 0 0 1560 870
use cc_inv_dco  cc_inv_dco_2
timestamp 1730452893
transform 1 0 3120 0 1 90
box 0 0 1560 870
use cc_inv_dco  cc_inv_dco_3
timestamp 1730452893
transform -1 0 3005 0 -1 -270
box 0 0 1560 870
use cc_inv_dco  cc_inv_dco_4
timestamp 1730452893
transform -1 0 4565 0 -1 -270
box 0 0 1560 870
<< labels >>
rlabel metal1 1405 -480 1405 -480 1 pn[4]
port 5 n
rlabel metal1 1400 -850 1400 -850 1 p[4]
port 10 n
rlabel metal1 4740 960 4740 960 1 VDDA
port 11 n
rlabel locali 1505 -100 1505 -100 3 VGND
port 12 e
<< end >>
