magic
tech sky130A
magscale 1 2
timestamp 1731569169
<< nwell >>
rect 3080 3700 3260 3820
rect 3080 3500 3256 3700
rect 7210 820 7340 1140
<< pwell >>
rect 3156 3390 3290 3394
rect 3100 3260 3290 3390
rect 3156 3258 3290 3260
rect 7170 580 7340 760
<< psubdiff >>
rect 3140 3342 3210 3380
rect 3140 3308 3164 3342
rect 3200 3308 3210 3342
rect 3140 3280 3210 3308
rect 3148 3276 3210 3280
rect 7230 690 7290 720
rect 7230 650 7240 690
rect 7280 650 7290 690
rect 7230 620 7290 650
<< nsubdiff >>
rect 3140 3662 3200 3696
rect 3140 3628 3154 3662
rect 3188 3628 3200 3662
rect 3140 3596 3200 3628
rect 7230 940 7290 970
rect 7230 900 7240 940
rect 7280 900 7290 940
rect 7230 870 7290 900
<< psubdiffcont >>
rect 3164 3308 3200 3342
rect 7240 650 7280 690
<< nsubdiffcont >>
rect 3154 3628 3188 3662
rect 7240 900 7280 940
<< locali >>
rect 3140 3670 3200 3696
rect 3730 3670 4190 3730
rect 3140 3630 3150 3670
rect 3190 3630 3200 3670
rect 3140 3628 3154 3630
rect 3188 3628 3200 3630
rect 3140 3596 3200 3628
rect 3690 3490 3760 3500
rect 3690 3450 3700 3490
rect 3740 3450 3760 3490
rect 3690 3440 3760 3450
rect 3140 3342 3210 3380
rect 3140 3308 3164 3342
rect 3200 3308 3210 3342
rect 3140 3270 3210 3308
rect 4130 3100 4190 3670
rect 10750 3520 13410 3540
rect 10750 3460 13210 3520
rect 13270 3460 13330 3520
rect 13390 3460 13410 3520
rect 10750 3440 13410 3460
rect 13310 3400 13410 3440
rect 13310 3340 13330 3400
rect 13390 3340 13410 3400
rect 13310 3320 13410 3340
rect 4120 3080 4200 3100
rect 4120 3040 4140 3080
rect 4180 3040 4200 3080
rect 4120 3020 4200 3040
rect 5980 -530 6080 1830
rect 7960 1370 8050 1390
rect 7960 1310 7970 1370
rect 8030 1310 8050 1370
rect 7960 1110 8050 1310
rect 7150 1040 8050 1110
rect 7230 940 7290 1040
rect 7230 900 7240 940
rect 7280 900 7290 940
rect 7230 870 7290 900
rect 7230 690 7290 720
rect 7230 650 7240 690
rect 7280 650 7290 690
rect 7230 620 7290 650
rect 7970 250 8050 1040
rect 6730 -190 6830 -170
rect 6730 -230 6760 -190
rect 6800 -230 6830 -190
rect 6730 -270 6830 -230
rect 7160 -490 7260 -470
rect 7160 -550 7180 -490
rect 7240 -550 7260 -490
rect 7160 -590 7260 -550
rect 7160 -610 7380 -590
rect 7160 -670 7180 -610
rect 7240 -670 7300 -610
rect 7360 -670 7380 -610
rect 7160 -690 7380 -670
rect 7160 -2080 7260 -690
rect 7160 -2100 7380 -2080
rect 7160 -2160 7180 -2100
rect 7240 -2160 7300 -2100
rect 7360 -2160 7380 -2100
rect 7160 -2180 7380 -2160
rect 7160 -2220 7260 -2180
rect 7160 -2280 7180 -2220
rect 7240 -2280 7260 -2220
rect 7160 -2300 7260 -2280
rect 6730 -2360 6830 -2340
rect 6730 -2400 6760 -2360
rect 6800 -2400 6830 -2360
rect 6730 -2410 6830 -2400
rect 6730 -2520 6830 -2510
rect 6730 -2560 6760 -2520
rect 6800 -2560 6830 -2520
rect 6730 -2580 6830 -2560
<< viali >>
rect 3150 3662 3190 3670
rect 3150 3630 3154 3662
rect 3154 3630 3188 3662
rect 3188 3630 3190 3662
rect 3330 3460 3370 3500
rect 3700 3450 3740 3490
rect 3164 3308 3200 3342
rect 4630 3560 4680 3610
rect 4630 3460 4680 3510
rect 4730 3460 4780 3510
rect 13210 3460 13270 3520
rect 13330 3460 13390 3520
rect 13330 3340 13390 3400
rect 4140 3040 4180 3080
rect 7970 1310 8030 1370
rect 7028 970 7062 1004
rect 7028 894 7062 928
rect 7240 900 7280 940
rect 6846 774 6880 808
rect 7240 650 7280 690
rect 6860 -140 6900 -100
rect 6760 -230 6800 -190
rect 7180 -550 7240 -490
rect 7180 -670 7240 -610
rect 7300 -670 7360 -610
rect 7180 -2160 7240 -2100
rect 7300 -2160 7360 -2100
rect 7180 -2280 7240 -2220
rect 6760 -2400 6800 -2360
rect 6760 -2560 6800 -2520
<< metal1 >>
rect 2220 3810 3300 3830
rect 2220 3750 2240 3810
rect 2300 3750 3300 3810
rect 2220 3740 3300 3750
rect 3740 3740 3920 3830
rect 3140 3670 3200 3740
rect 3140 3630 3150 3670
rect 3190 3630 3200 3670
rect 3140 3596 3200 3630
rect 3300 3500 3400 3540
rect 3850 3500 3920 3740
rect 4610 3610 4690 3630
rect 4610 3560 4630 3610
rect 4680 3560 4690 3610
rect 4610 3520 4690 3560
rect 13190 3520 13410 3540
rect 3300 3490 3330 3500
rect 2890 3460 3330 3490
rect 3370 3460 3400 3500
rect 2890 3430 3400 3460
rect 3680 3490 3920 3500
rect 3680 3450 3700 3490
rect 3740 3450 3920 3490
rect 3680 3430 3920 3450
rect 4320 3510 4800 3520
rect 4320 3460 4630 3510
rect 4680 3460 4730 3510
rect 4780 3460 4800 3510
rect 4320 3440 4800 3460
rect 13190 3460 13210 3520
rect 13270 3460 13330 3520
rect 13390 3460 13410 3520
rect 13190 3440 13410 3460
rect 3140 3342 3210 3380
rect 3140 3308 3164 3342
rect 3200 3308 3210 3342
rect 3140 3280 3210 3308
rect 4320 3280 4420 3440
rect 3100 3190 3300 3280
rect 3740 3190 4420 3280
rect 13310 3400 13410 3440
rect 13310 3340 13330 3400
rect 13390 3340 13410 3400
rect 4220 1120 4300 2280
rect 7840 1370 8050 1390
rect 7840 1310 7970 1370
rect 8030 1310 8050 1370
rect 7840 1300 8050 1310
rect 4220 1040 6490 1120
rect 6410 830 6490 1040
rect 7020 1004 7070 1020
rect 7020 970 7028 1004
rect 7062 970 7070 1004
rect 7020 928 7070 970
rect 7020 894 7028 928
rect 7062 894 7070 928
rect 6410 828 6830 830
rect 6410 808 6896 828
rect 6410 774 6846 808
rect 6880 774 6896 808
rect 7020 820 7070 894
rect 7230 940 7290 970
rect 7230 900 7240 940
rect 7280 900 7290 940
rect 7230 870 7290 900
rect 7350 820 8270 850
rect 7020 780 8270 820
rect 7037 778 8270 780
rect 6410 756 6896 774
rect 6410 750 6830 756
rect 7350 750 8270 778
rect 7230 690 7290 720
rect 2850 590 5590 690
rect 7230 650 7240 690
rect 7280 650 7290 690
rect 7230 600 7290 650
rect 2230 290 2240 350
rect 2300 290 2310 350
rect 2850 160 2950 590
rect 2640 60 2950 160
rect 3750 60 4390 160
rect 5490 150 5590 590
rect 6730 -70 6830 600
rect 7170 510 7290 600
rect 8170 10 8270 750
rect 6830 -100 6930 -70
rect 6830 -140 6860 -100
rect 6900 -140 6930 -100
rect 6830 -170 6930 -140
rect 11500 -390 11600 -370
rect 11500 -450 11520 -390
rect 11580 -450 11600 -390
rect 11500 -470 11600 -450
rect 1240 -1880 1320 -1720
rect 6730 -2360 6830 -772
rect 8150 -1440 8250 -1420
rect 8150 -1500 8170 -1440
rect 8230 -1500 8250 -1440
rect 8150 -2340 8250 -1500
rect 6730 -2400 6760 -2360
rect 6800 -2400 6830 -2360
rect 6730 -2520 6830 -2400
rect 6730 -2534 6760 -2520
rect 6800 -2534 6830 -2520
rect 11500 -2820 11600 -2740
rect 2800 -4370 2900 -3510
rect 6730 -4370 6830 -3180
rect 13310 -4370 13410 3340
rect 2800 -4470 13410 -4370
<< via1 >>
rect 2240 3750 2300 3810
rect 7970 1310 8030 1370
rect 2240 290 2300 350
rect 11520 -450 11580 -390
rect 8170 -1500 8230 -1440
<< metal2 >>
rect 2220 3810 2320 3830
rect 2220 3750 2240 3810
rect 2300 3750 2320 3810
rect 2220 1390 2320 3750
rect 2220 1370 8050 1390
rect 2220 1310 7970 1370
rect 8030 1310 8050 1370
rect 2220 1300 8050 1310
rect 2220 350 2320 1300
rect 2220 290 2240 350
rect 2300 290 2320 350
rect 2220 280 2320 290
rect 11500 -390 12010 -370
rect 11500 -450 11520 -390
rect 11580 -450 12010 -390
rect 11500 -470 12010 -450
rect 11910 -1420 12010 -470
rect 8150 -1440 12010 -1420
rect 8150 -1500 8170 -1440
rect 8230 -1500 12010 -1440
rect 8150 -1520 12010 -1500
use ALib_IDAC  ALib_IDAC_0
timestamp 1731569169
transform 1 0 2860 0 1 -380
box -1860 -3160 3220 740
use DLib_freqDiv2  DLib_freqDiv2_0
timestamp 1731569169
transform 1 0 8320 0 1 -2610
box -1590 -1450 4400 640
use DLib_freqDiv2  DLib_freqDiv2_1
timestamp 1731569169
transform 1 0 8320 0 1 -270
box -1590 -1450 4400 640
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6808 0 1 558
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  sky130_fd_sc_hd__einvp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3288 0 1 3238
box -38 -48 498 592
use x5s_cc_osc_dco  x5s_cc_osc_dco_0
timestamp 1731473513
transform 1 0 1680 0 1 4060
box -500 -2280 10480 1920
<< labels >>
rlabel metal1 2950 690 2950 690 1 Vbs_12
port 1 n
rlabel metal1 4030 160 4030 160 1 Vbs_34
port 2 n
rlabel metal1 1240 -1750 1240 -1750 7 Dctrl
port 4 w
rlabel metal1 2930 3490 2930 3490 1 ENB
port 5 n
rlabel metal1 3880 3830 3880 3830 1 VDDA
port 6 n
rlabel metal1 2940 -4370 2940 -4370 1 GND
port 7 n
rlabel metal1 11580 -2740 11580 -2740 1 pha_DCO
port 3 n
<< end >>
