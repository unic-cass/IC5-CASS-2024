magic
tech sky130A
timestamp 1730442115
<< nwell >>
rect -130 -45 425 535
<< pwell >>
rect -130 -550 425 -70
<< nmos >>
rect 0 -510 365 -110
<< pmos >>
rect 0 -5 365 495
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -320 0 -300
rect -40 -340 -30 -320
rect -10 -340 0 -320
rect -40 -360 0 -340
rect -40 -380 -30 -360
rect -10 -380 0 -360
rect -40 -400 0 -380
rect -40 -420 -30 -400
rect -10 -420 0 -400
rect -40 -440 0 -420
rect -40 -460 -30 -440
rect -10 -460 0 -440
rect -40 -480 0 -460
rect -40 -500 -30 -480
rect -10 -500 0 -480
rect -40 -510 0 -500
rect 365 -120 405 -110
rect 365 -140 375 -120
rect 395 -140 405 -120
rect 365 -160 405 -140
rect 365 -180 375 -160
rect 395 -180 405 -160
rect 365 -200 405 -180
rect 365 -220 375 -200
rect 395 -220 405 -200
rect 365 -240 405 -220
rect 365 -260 375 -240
rect 395 -260 405 -240
rect 365 -280 405 -260
rect 365 -300 375 -280
rect 395 -300 405 -280
rect 365 -320 405 -300
rect 365 -340 375 -320
rect 395 -340 405 -320
rect 365 -360 405 -340
rect 365 -380 375 -360
rect 395 -380 405 -360
rect 365 -400 405 -380
rect 365 -420 375 -400
rect 395 -420 405 -400
rect 365 -440 405 -420
rect 365 -460 375 -440
rect 395 -460 405 -440
rect 365 -480 405 -460
rect 365 -500 375 -480
rect 395 -500 405 -480
rect 365 -510 405 -500
<< pdiff >>
rect -40 485 0 495
rect -40 465 -30 485
rect -10 465 0 485
rect -40 445 0 465
rect -40 425 -30 445
rect -10 425 0 445
rect -40 405 0 425
rect -40 385 -30 405
rect -10 385 0 405
rect -40 365 0 385
rect -40 345 -30 365
rect -10 345 0 365
rect -40 325 0 345
rect -40 305 -30 325
rect -10 305 0 325
rect -40 285 0 305
rect -40 265 -30 285
rect -10 265 0 285
rect -40 245 0 265
rect -40 225 -30 245
rect -10 225 0 245
rect -40 205 0 225
rect -40 185 -30 205
rect -10 185 0 205
rect -40 165 0 185
rect -40 145 -30 165
rect -10 145 0 165
rect -40 125 0 145
rect -40 105 -30 125
rect -10 105 0 125
rect -40 85 0 105
rect -40 65 -30 85
rect -10 65 0 85
rect -40 45 0 65
rect -40 25 -30 45
rect -10 25 0 45
rect -40 -5 0 25
rect 365 485 405 495
rect 365 465 375 485
rect 395 465 405 485
rect 365 445 405 465
rect 365 425 375 445
rect 395 425 405 445
rect 365 405 405 425
rect 365 385 375 405
rect 395 385 405 405
rect 365 365 405 385
rect 365 345 375 365
rect 395 345 405 365
rect 365 325 405 345
rect 365 305 375 325
rect 395 305 405 325
rect 365 285 405 305
rect 365 265 375 285
rect 395 265 405 285
rect 365 245 405 265
rect 365 225 375 245
rect 395 225 405 245
rect 365 205 405 225
rect 365 185 375 205
rect 395 185 405 205
rect 365 165 405 185
rect 365 145 375 165
rect 395 145 405 165
rect 365 125 405 145
rect 365 105 375 125
rect 395 105 405 125
rect 365 85 405 105
rect 365 65 375 85
rect 395 65 405 85
rect 365 45 405 65
rect 365 25 375 45
rect 395 25 405 45
rect 365 -5 405 25
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect -30 -340 -10 -320
rect -30 -380 -10 -360
rect -30 -420 -10 -400
rect -30 -460 -10 -440
rect -30 -500 -10 -480
rect 375 -140 395 -120
rect 375 -180 395 -160
rect 375 -220 395 -200
rect 375 -260 395 -240
rect 375 -300 395 -280
rect 375 -340 395 -320
rect 375 -380 395 -360
rect 375 -420 395 -400
rect 375 -460 395 -440
rect 375 -500 395 -480
<< pdiffc >>
rect -30 465 -10 485
rect -30 425 -10 445
rect -30 385 -10 405
rect -30 345 -10 365
rect -30 305 -10 325
rect -30 265 -10 285
rect -30 225 -10 245
rect -30 185 -10 205
rect -30 145 -10 165
rect -30 105 -10 125
rect -30 65 -10 85
rect -30 25 -10 45
rect 375 465 395 485
rect 375 425 395 445
rect 375 385 395 405
rect 375 345 395 365
rect 375 305 395 325
rect 375 265 395 285
rect 375 225 395 245
rect 375 185 395 205
rect 375 145 395 165
rect 375 105 395 125
rect 375 65 395 85
rect 375 25 395 45
<< psubdiff >>
rect -110 -480 -70 -465
rect -110 -500 -100 -480
rect -80 -500 -70 -480
rect -110 -515 -70 -500
<< nsubdiff >>
rect -110 485 -70 500
rect -110 465 -100 485
rect -80 465 -70 485
rect -110 450 -70 465
<< psubdiffcont >>
rect -100 -500 -80 -480
<< nsubdiffcont >>
rect -100 465 -80 485
<< poly >>
rect 0 495 365 535
rect 0 -110 365 -5
rect 0 -550 365 -510
<< locali >>
rect -110 495 -70 500
rect -110 485 0 495
rect -110 465 -100 485
rect -80 465 -30 485
rect -10 465 0 485
rect -110 450 0 465
rect -40 445 0 450
rect -40 425 -30 445
rect -10 425 0 445
rect -40 405 0 425
rect -40 385 -30 405
rect -10 385 0 405
rect -40 365 0 385
rect -40 345 -30 365
rect -10 345 0 365
rect -40 325 0 345
rect -40 305 -30 325
rect -10 305 0 325
rect -40 285 0 305
rect -40 265 -30 285
rect -10 265 0 285
rect -40 245 0 265
rect -40 225 -30 245
rect -10 225 0 245
rect -40 205 0 225
rect -40 185 -30 205
rect -10 185 0 205
rect -40 165 0 185
rect -40 145 -30 165
rect -10 145 0 165
rect -40 125 0 145
rect -40 105 -30 125
rect -10 105 0 125
rect -40 85 0 105
rect -40 65 -30 85
rect -10 65 0 85
rect -40 45 0 65
rect -40 25 -30 45
rect -10 25 0 45
rect -40 -5 0 25
rect 365 485 405 495
rect 365 465 375 485
rect 395 465 405 485
rect 365 445 405 465
rect 365 425 375 445
rect 395 425 405 445
rect 365 405 405 425
rect 365 385 375 405
rect 395 385 405 405
rect 365 365 405 385
rect 365 345 375 365
rect 395 345 405 365
rect 365 325 405 345
rect 365 305 375 325
rect 395 305 405 325
rect 365 285 405 305
rect 365 265 375 285
rect 395 265 405 285
rect 365 245 405 265
rect 365 225 375 245
rect 395 225 405 245
rect 365 205 405 225
rect 365 185 375 205
rect 395 185 405 205
rect 365 165 405 185
rect 365 145 375 165
rect 395 145 405 165
rect 365 125 405 145
rect 365 105 375 125
rect 395 105 405 125
rect 365 85 405 105
rect 365 65 375 85
rect 395 65 405 85
rect 365 45 405 65
rect 365 25 375 45
rect 395 25 405 45
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -320 0 -300
rect -40 -340 -30 -320
rect -10 -340 0 -320
rect -40 -360 0 -340
rect -40 -380 -30 -360
rect -10 -380 0 -360
rect -40 -400 0 -380
rect -40 -420 -30 -400
rect -10 -420 0 -400
rect -40 -440 0 -420
rect -40 -460 -30 -440
rect -10 -460 0 -440
rect -110 -480 -70 -465
rect -110 -500 -100 -480
rect -80 -500 -70 -480
rect -110 -515 -70 -500
rect -40 -480 0 -460
rect -40 -500 -30 -480
rect -10 -500 0 -480
rect -40 -510 0 -500
rect 365 -120 405 25
rect 365 -140 375 -120
rect 395 -140 405 -120
rect 365 -160 405 -140
rect 365 -180 375 -160
rect 395 -180 405 -160
rect 365 -200 405 -180
rect 365 -220 375 -200
rect 395 -220 405 -200
rect 365 -240 405 -220
rect 365 -260 375 -240
rect 395 -260 405 -240
rect 365 -280 405 -260
rect 365 -300 375 -280
rect 395 -300 405 -280
rect 365 -320 405 -300
rect 365 -340 375 -320
rect 395 -340 405 -320
rect 365 -360 405 -340
rect 365 -380 375 -360
rect 395 -380 405 -360
rect 365 -400 405 -380
rect 365 -420 375 -400
rect 395 -420 405 -400
rect 365 -440 405 -420
rect 365 -460 375 -440
rect 395 -460 405 -440
rect 365 -480 405 -460
rect 365 -500 375 -480
rect 395 -500 405 -480
rect 365 -510 405 -500
<< viali >>
rect -100 465 -80 485
rect -100 -500 -80 -480
<< metal1 >>
rect -110 485 -70 500
rect -110 465 -100 485
rect -80 465 -70 485
rect -110 450 -70 465
rect -110 -480 -70 -465
rect -110 -500 -100 -480
rect -80 -500 -70 -480
rect -110 -515 -70 -500
<< labels >>
rlabel poly 0 -55 0 -55 7 A
port 1 w
rlabel locali 405 -60 405 -60 3 Y
port 2 e
rlabel locali -20 -510 -20 -510 5 VGND
port 3 s
rlabel metal1 -90 500 -90 500 1 VDDA
port 4 n
rlabel metal1 -90 -515 -90 -515 5 GND
port 5 s
<< end >>
