magic
tech sky130A
magscale 1 2
timestamp 1731481839
<< obsli1 >>
rect 1104 2159 254840 255697
<< obsm1 >>
rect 1104 1368 254840 256012
<< metal2 >>
rect 63958 257378 64014 258178
rect 191930 257378 191986 258178
rect 2410 0 2466 800
rect 4802 0 4858 800
rect 7194 0 7250 800
rect 9586 0 9642 800
rect 11978 0 12034 800
rect 14370 0 14426 800
rect 16762 0 16818 800
rect 19154 0 19210 800
rect 21546 0 21602 800
rect 23938 0 23994 800
rect 26330 0 26386 800
rect 28722 0 28778 800
rect 31114 0 31170 800
rect 33506 0 33562 800
rect 35898 0 35954 800
rect 38290 0 38346 800
rect 40682 0 40738 800
rect 43074 0 43130 800
rect 45466 0 45522 800
rect 47858 0 47914 800
rect 50250 0 50306 800
rect 52642 0 52698 800
rect 55034 0 55090 800
rect 57426 0 57482 800
rect 59818 0 59874 800
rect 62210 0 62266 800
rect 64602 0 64658 800
rect 66994 0 67050 800
rect 69386 0 69442 800
rect 71778 0 71834 800
rect 74170 0 74226 800
rect 76562 0 76618 800
rect 78954 0 79010 800
rect 81346 0 81402 800
rect 83738 0 83794 800
rect 86130 0 86186 800
rect 88522 0 88578 800
rect 90914 0 90970 800
rect 93306 0 93362 800
rect 95698 0 95754 800
rect 98090 0 98146 800
rect 100482 0 100538 800
rect 102874 0 102930 800
rect 105266 0 105322 800
rect 107658 0 107714 800
rect 110050 0 110106 800
rect 112442 0 112498 800
rect 114834 0 114890 800
rect 117226 0 117282 800
rect 119618 0 119674 800
rect 122010 0 122066 800
rect 124402 0 124458 800
rect 126794 0 126850 800
rect 129186 0 129242 800
rect 131578 0 131634 800
rect 133970 0 134026 800
rect 136362 0 136418 800
rect 138754 0 138810 800
rect 141146 0 141202 800
rect 143538 0 143594 800
rect 145930 0 145986 800
rect 148322 0 148378 800
rect 150714 0 150770 800
rect 153106 0 153162 800
rect 155498 0 155554 800
rect 157890 0 157946 800
rect 160282 0 160338 800
rect 162674 0 162730 800
rect 165066 0 165122 800
rect 167458 0 167514 800
rect 169850 0 169906 800
rect 172242 0 172298 800
rect 174634 0 174690 800
rect 177026 0 177082 800
rect 179418 0 179474 800
rect 181810 0 181866 800
rect 184202 0 184258 800
rect 186594 0 186650 800
rect 188986 0 189042 800
rect 191378 0 191434 800
rect 193770 0 193826 800
rect 196162 0 196218 800
rect 198554 0 198610 800
rect 200946 0 201002 800
rect 203338 0 203394 800
rect 205730 0 205786 800
rect 208122 0 208178 800
rect 210514 0 210570 800
rect 212906 0 212962 800
rect 215298 0 215354 800
rect 217690 0 217746 800
rect 220082 0 220138 800
rect 222474 0 222530 800
rect 224866 0 224922 800
rect 227258 0 227314 800
rect 229650 0 229706 800
rect 232042 0 232098 800
rect 234434 0 234490 800
rect 236826 0 236882 800
rect 239218 0 239274 800
rect 241610 0 241666 800
rect 244002 0 244058 800
rect 246394 0 246450 800
rect 248786 0 248842 800
rect 251178 0 251234 800
rect 253570 0 253626 800
<< obsm2 >>
rect 2410 257322 63902 257530
rect 64070 257322 191874 257530
rect 192042 257322 253624 257530
rect 2410 856 253624 257322
rect 2522 734 4746 856
rect 4914 734 7138 856
rect 7306 734 9530 856
rect 9698 734 11922 856
rect 12090 734 14314 856
rect 14482 734 16706 856
rect 16874 734 19098 856
rect 19266 734 21490 856
rect 21658 734 23882 856
rect 24050 734 26274 856
rect 26442 734 28666 856
rect 28834 734 31058 856
rect 31226 734 33450 856
rect 33618 734 35842 856
rect 36010 734 38234 856
rect 38402 734 40626 856
rect 40794 734 43018 856
rect 43186 734 45410 856
rect 45578 734 47802 856
rect 47970 734 50194 856
rect 50362 734 52586 856
rect 52754 734 54978 856
rect 55146 734 57370 856
rect 57538 734 59762 856
rect 59930 734 62154 856
rect 62322 734 64546 856
rect 64714 734 66938 856
rect 67106 734 69330 856
rect 69498 734 71722 856
rect 71890 734 74114 856
rect 74282 734 76506 856
rect 76674 734 78898 856
rect 79066 734 81290 856
rect 81458 734 83682 856
rect 83850 734 86074 856
rect 86242 734 88466 856
rect 88634 734 90858 856
rect 91026 734 93250 856
rect 93418 734 95642 856
rect 95810 734 98034 856
rect 98202 734 100426 856
rect 100594 734 102818 856
rect 102986 734 105210 856
rect 105378 734 107602 856
rect 107770 734 109994 856
rect 110162 734 112386 856
rect 112554 734 114778 856
rect 114946 734 117170 856
rect 117338 734 119562 856
rect 119730 734 121954 856
rect 122122 734 124346 856
rect 124514 734 126738 856
rect 126906 734 129130 856
rect 129298 734 131522 856
rect 131690 734 133914 856
rect 134082 734 136306 856
rect 136474 734 138698 856
rect 138866 734 141090 856
rect 141258 734 143482 856
rect 143650 734 145874 856
rect 146042 734 148266 856
rect 148434 734 150658 856
rect 150826 734 153050 856
rect 153218 734 155442 856
rect 155610 734 157834 856
rect 158002 734 160226 856
rect 160394 734 162618 856
rect 162786 734 165010 856
rect 165178 734 167402 856
rect 167570 734 169794 856
rect 169962 734 172186 856
rect 172354 734 174578 856
rect 174746 734 176970 856
rect 177138 734 179362 856
rect 179530 734 181754 856
rect 181922 734 184146 856
rect 184314 734 186538 856
rect 186706 734 188930 856
rect 189098 734 191322 856
rect 191490 734 193714 856
rect 193882 734 196106 856
rect 196274 734 198498 856
rect 198666 734 200890 856
rect 201058 734 203282 856
rect 203450 734 205674 856
rect 205842 734 208066 856
rect 208234 734 210458 856
rect 210626 734 212850 856
rect 213018 734 215242 856
rect 215410 734 217634 856
rect 217802 734 220026 856
rect 220194 734 222418 856
rect 222586 734 224810 856
rect 224978 734 227202 856
rect 227370 734 229594 856
rect 229762 734 231986 856
rect 232154 734 234378 856
rect 234546 734 236770 856
rect 236938 734 239162 856
rect 239330 734 241554 856
rect 241722 734 243946 856
rect 244114 734 246338 856
rect 246506 734 248730 856
rect 248898 734 251122 856
rect 251290 734 253514 856
<< metal3 >>
rect 0 128936 800 129056
<< obsm3 >>
rect 800 129136 252527 255713
rect 880 128856 252527 129136
rect 800 1803 252527 128856
<< metal4 >>
rect 4208 2128 4528 255728
rect 19568 2128 19888 255728
rect 34928 2128 35248 255728
rect 50288 2128 50608 255728
rect 65648 2128 65968 255728
rect 81008 2128 81328 255728
rect 96368 2128 96688 255728
rect 111728 2128 112048 255728
rect 127088 2128 127408 255728
rect 142448 2128 142768 255728
rect 157808 2128 158128 255728
rect 173168 2128 173488 255728
rect 188528 2128 188848 255728
rect 203888 2128 204208 255728
rect 219248 2128 219568 255728
rect 234608 2128 234928 255728
rect 249968 2128 250288 255728
<< obsm4 >>
rect 9443 2891 19488 255373
rect 19968 2891 34848 255373
rect 35328 2891 50208 255373
rect 50688 2891 65568 255373
rect 66048 2891 80928 255373
rect 81408 2891 96288 255373
rect 96768 2891 111648 255373
rect 112128 2891 127008 255373
rect 127488 2891 142368 255373
rect 142848 2891 157728 255373
rect 158208 2891 173088 255373
rect 173568 2891 188448 255373
rect 188928 2891 203808 255373
rect 204288 2891 219168 255373
rect 219648 2891 234528 255373
rect 235008 2891 248709 255373
<< labels >>
rlabel metal2 s 63958 257378 64014 258178 6 phase_in
port 1 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 user_clock2
port 2 nsew signal input
rlabel metal4 s 4208 2128 4528 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 255728 6 vccd1
port 3 nsew power bidirectional
rlabel metal2 s 191930 257378 191986 258178 6 vco_enb_o
port 4 nsew signal output
rlabel metal4 s 19568 2128 19888 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 255728 6 vssd1
port 5 nsew ground bidirectional
rlabel metal2 s 2410 0 2466 800 6 wb_clk_i
port 6 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wb_rst_i
port 7 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_ack_o
port 8 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[0]
port 9 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 wbs_adr_i[10]
port 10 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 wbs_adr_i[11]
port 11 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 wbs_adr_i[12]
port 12 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 wbs_adr_i[13]
port 13 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 wbs_adr_i[14]
port 14 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 wbs_adr_i[15]
port 15 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 wbs_adr_i[16]
port 16 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 wbs_adr_i[17]
port 17 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 wbs_adr_i[18]
port 18 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 wbs_adr_i[19]
port 19 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[1]
port 20 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 wbs_adr_i[20]
port 21 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 wbs_adr_i[21]
port 22 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 wbs_adr_i[22]
port 23 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 wbs_adr_i[23]
port 24 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 wbs_adr_i[24]
port 25 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 wbs_adr_i[25]
port 26 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 wbs_adr_i[26]
port 27 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 wbs_adr_i[27]
port 28 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 wbs_adr_i[28]
port 29 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 wbs_adr_i[29]
port 30 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[2]
port 31 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 wbs_adr_i[30]
port 32 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 wbs_adr_i[31]
port 33 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_adr_i[3]
port 34 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_adr_i[4]
port 35 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 wbs_adr_i[5]
port 36 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_adr_i[6]
port 37 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 wbs_adr_i[7]
port 38 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 wbs_adr_i[8]
port 39 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 wbs_adr_i[9]
port 40 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_cyc_i
port 41 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[0]
port 42 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_dat_i[10]
port 43 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 wbs_dat_i[11]
port 44 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 wbs_dat_i[12]
port 45 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 wbs_dat_i[13]
port 46 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 wbs_dat_i[14]
port 47 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 wbs_dat_i[15]
port 48 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 wbs_dat_i[16]
port 49 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 wbs_dat_i[17]
port 50 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 wbs_dat_i[18]
port 51 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 wbs_dat_i[19]
port 52 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[1]
port 53 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 wbs_dat_i[20]
port 54 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 wbs_dat_i[21]
port 55 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 wbs_dat_i[22]
port 56 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 wbs_dat_i[23]
port 57 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 wbs_dat_i[24]
port 58 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 wbs_dat_i[25]
port 59 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 wbs_dat_i[26]
port 60 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 wbs_dat_i[27]
port 61 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 wbs_dat_i[28]
port 62 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 wbs_dat_i[29]
port 63 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[2]
port 64 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 wbs_dat_i[30]
port 65 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 wbs_dat_i[31]
port 66 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[3]
port 67 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_i[4]
port 68 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_i[5]
port 69 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_i[6]
port 70 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_dat_i[7]
port 71 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 wbs_dat_i[8]
port 72 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_i[9]
port 73 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[0]
port 74 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 wbs_dat_o[10]
port 75 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 wbs_dat_o[11]
port 76 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 wbs_dat_o[12]
port 77 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 wbs_dat_o[13]
port 78 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_o[14]
port 79 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 wbs_dat_o[15]
port 80 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 wbs_dat_o[16]
port 81 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 wbs_dat_o[17]
port 82 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 wbs_dat_o[18]
port 83 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 wbs_dat_o[19]
port 84 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[1]
port 85 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 wbs_dat_o[20]
port 86 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 wbs_dat_o[21]
port 87 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 wbs_dat_o[22]
port 88 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 wbs_dat_o[23]
port 89 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 wbs_dat_o[24]
port 90 nsew signal output
rlabel metal2 s 210514 0 210570 800 6 wbs_dat_o[25]
port 91 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 wbs_dat_o[26]
port 92 nsew signal output
rlabel metal2 s 224866 0 224922 800 6 wbs_dat_o[27]
port 93 nsew signal output
rlabel metal2 s 232042 0 232098 800 6 wbs_dat_o[28]
port 94 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 wbs_dat_o[29]
port 95 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[2]
port 96 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 wbs_dat_o[30]
port 97 nsew signal output
rlabel metal2 s 253570 0 253626 800 6 wbs_dat_o[31]
port 98 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_o[3]
port 99 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_o[4]
port 100 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 wbs_dat_o[5]
port 101 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 wbs_dat_o[6]
port 102 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 wbs_dat_o[7]
port 103 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_o[8]
port 104 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[9]
port 105 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_sel_i[0]
port 106 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_sel_i[1]
port 107 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_sel_i[2]
port 108 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_sel_i[3]
port 109 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_stb_i
port 110 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_we_i
port 111 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 256034 258178
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 191870910
string GDS_FILE /home/admin/projects/IC5-CASS-2024/openlane/vco_adc_wrapper/runs/24_11_13_11_29/results/signoff/vco_adc_wrapper.magic.gds
string GDS_START 1248028
<< end >>

