magic
tech sky130A
magscale 1 2
timestamp 1731299803
<< nwell >>
rect 1066 132997 133070 133563
rect 1066 131909 133070 132475
rect 1066 130821 133070 131387
rect 1066 129733 133070 130299
rect 1066 128645 133070 129211
rect 1066 127557 133070 128123
rect 1066 126469 133070 127035
rect 1066 125381 133070 125947
rect 1066 124293 133070 124859
rect 1066 123205 133070 123771
rect 1066 122117 133070 122683
rect 1066 121029 133070 121595
rect 1066 119941 133070 120507
rect 1066 118853 133070 119419
rect 1066 117765 133070 118331
rect 1066 116677 133070 117243
rect 1066 115589 133070 116155
rect 1066 114501 133070 115067
rect 1066 113413 133070 113979
rect 1066 112325 133070 112891
rect 1066 111237 133070 111803
rect 1066 110149 133070 110715
rect 1066 109061 133070 109627
rect 1066 107973 133070 108539
rect 1066 106885 133070 107451
rect 1066 105797 133070 106363
rect 1066 104709 133070 105275
rect 1066 103621 133070 104187
rect 1066 102533 133070 103099
rect 1066 101445 133070 102011
rect 1066 100357 133070 100923
rect 1066 99269 133070 99835
rect 1066 98181 133070 98747
rect 1066 97093 133070 97659
rect 1066 96005 133070 96571
rect 1066 94917 133070 95483
rect 1066 93829 133070 94395
rect 1066 92741 133070 93307
rect 1066 91653 133070 92219
rect 1066 90565 133070 91131
rect 1066 89477 133070 90043
rect 1066 88389 133070 88955
rect 1066 87301 133070 87867
rect 1066 86213 133070 86779
rect 1066 85125 133070 85691
rect 1066 84037 133070 84603
rect 1066 82949 133070 83515
rect 1066 81861 133070 82427
rect 1066 80773 133070 81339
rect 1066 79685 133070 80251
rect 1066 78597 133070 79163
rect 1066 77509 133070 78075
rect 1066 76421 133070 76987
rect 1066 75333 133070 75899
rect 1066 74245 133070 74811
rect 1066 73157 133070 73723
rect 1066 72069 133070 72635
rect 1066 70981 133070 71547
rect 1066 69893 133070 70459
rect 1066 68805 133070 69371
rect 1066 67717 133070 68283
rect 1066 66629 133070 67195
rect 1066 65541 133070 66107
rect 1066 64453 133070 65019
rect 1066 63365 133070 63931
rect 1066 62277 133070 62843
rect 1066 61189 133070 61755
rect 1066 60101 133070 60667
rect 1066 59013 133070 59579
rect 1066 57925 133070 58491
rect 1066 56837 133070 57403
rect 1066 55749 133070 56315
rect 1066 54661 133070 55227
rect 1066 53573 133070 54139
rect 1066 52485 133070 53051
rect 1066 51397 133070 51963
rect 1066 50309 133070 50875
rect 1066 49221 133070 49787
rect 1066 48133 133070 48699
rect 1066 47045 133070 47611
rect 1066 45957 133070 46523
rect 1066 44869 133070 45435
rect 1066 43781 133070 44347
rect 1066 42693 133070 43259
rect 1066 41605 133070 42171
rect 1066 40517 133070 41083
rect 1066 39429 133070 39995
rect 1066 38341 133070 38907
rect 1066 37253 133070 37819
rect 1066 36165 133070 36731
rect 1066 35077 133070 35643
rect 1066 33989 133070 34555
rect 1066 32901 133070 33467
rect 1066 31813 133070 32379
rect 1066 30725 133070 31291
rect 1066 29637 133070 30203
rect 1066 28549 133070 29115
rect 1066 27461 133070 28027
rect 1066 26373 133070 26939
rect 1066 25285 133070 25851
rect 1066 24197 133070 24763
rect 1066 23109 133070 23675
rect 1066 22021 133070 22587
rect 1066 20933 133070 21499
rect 1066 19845 133070 20411
rect 1066 18757 133070 19323
rect 1066 17669 133070 18235
rect 1066 16581 133070 17147
rect 1066 15493 133070 16059
rect 1066 14405 133070 14971
rect 1066 13317 133070 13883
rect 1066 12229 133070 12795
rect 1066 11141 133070 11707
rect 1066 10053 133070 10619
rect 1066 8965 133070 9531
rect 1066 7877 133070 8443
rect 1066 6789 133070 7355
rect 1066 5701 133070 6267
rect 1066 4613 133070 5179
rect 1066 3525 133070 4091
rect 1066 2437 133070 3003
<< obsli1 >>
rect 1104 2159 133032 133841
<< obsm1 >>
rect 1104 1776 133032 133872
<< metal2 >>
rect 2410 135512 2466 136312
rect 4066 135512 4122 136312
rect 5722 135512 5778 136312
rect 7378 135512 7434 136312
rect 9034 135512 9090 136312
rect 10690 135512 10746 136312
rect 12346 135512 12402 136312
rect 14002 135512 14058 136312
rect 15658 135512 15714 136312
rect 17314 135512 17370 136312
rect 18970 135512 19026 136312
rect 20626 135512 20682 136312
rect 22282 135512 22338 136312
rect 23938 135512 23994 136312
rect 25594 135512 25650 136312
rect 27250 135512 27306 136312
rect 28906 135512 28962 136312
rect 30562 135512 30618 136312
rect 32218 135512 32274 136312
rect 33874 135512 33930 136312
rect 35530 135512 35586 136312
rect 37186 135512 37242 136312
rect 38842 135512 38898 136312
rect 40498 135512 40554 136312
rect 42154 135512 42210 136312
rect 43810 135512 43866 136312
rect 45466 135512 45522 136312
rect 47122 135512 47178 136312
rect 48778 135512 48834 136312
rect 50434 135512 50490 136312
rect 52090 135512 52146 136312
rect 53746 135512 53802 136312
rect 55402 135512 55458 136312
rect 57058 135512 57114 136312
rect 58714 135512 58770 136312
rect 60370 135512 60426 136312
rect 62026 135512 62082 136312
rect 63682 135512 63738 136312
rect 65338 135512 65394 136312
rect 66994 135512 67050 136312
rect 68650 135512 68706 136312
rect 70306 135512 70362 136312
rect 71962 135512 72018 136312
rect 73618 135512 73674 136312
rect 75274 135512 75330 136312
rect 76930 135512 76986 136312
rect 78586 135512 78642 136312
rect 80242 135512 80298 136312
rect 81898 135512 81954 136312
rect 83554 135512 83610 136312
rect 85210 135512 85266 136312
rect 86866 135512 86922 136312
rect 88522 135512 88578 136312
rect 90178 135512 90234 136312
rect 91834 135512 91890 136312
rect 93490 135512 93546 136312
rect 95146 135512 95202 136312
rect 96802 135512 96858 136312
rect 98458 135512 98514 136312
rect 100114 135512 100170 136312
rect 101770 135512 101826 136312
rect 103426 135512 103482 136312
rect 105082 135512 105138 136312
rect 106738 135512 106794 136312
rect 108394 135512 108450 136312
rect 110050 135512 110106 136312
rect 111706 135512 111762 136312
rect 113362 135512 113418 136312
rect 115018 135512 115074 136312
rect 116674 135512 116730 136312
rect 118330 135512 118386 136312
rect 119986 135512 120042 136312
rect 121642 135512 121698 136312
rect 123298 135512 123354 136312
rect 124954 135512 125010 136312
rect 126610 135512 126666 136312
rect 128266 135512 128322 136312
rect 129922 135512 129978 136312
rect 131578 135512 131634 136312
rect 1214 0 1270 800
rect 3238 0 3294 800
rect 5262 0 5318 800
rect 7286 0 7342 800
rect 9310 0 9366 800
rect 11334 0 11390 800
rect 13358 0 13414 800
rect 15382 0 15438 800
rect 17406 0 17462 800
rect 19430 0 19486 800
rect 21454 0 21510 800
rect 23478 0 23534 800
rect 25502 0 25558 800
rect 27526 0 27582 800
rect 29550 0 29606 800
rect 31574 0 31630 800
rect 33598 0 33654 800
rect 35622 0 35678 800
rect 37646 0 37702 800
rect 39670 0 39726 800
rect 41694 0 41750 800
rect 43718 0 43774 800
rect 45742 0 45798 800
rect 47766 0 47822 800
rect 49790 0 49846 800
rect 51814 0 51870 800
rect 53838 0 53894 800
rect 55862 0 55918 800
rect 57886 0 57942 800
rect 59910 0 59966 800
rect 61934 0 61990 800
rect 63958 0 64014 800
rect 65982 0 66038 800
rect 68006 0 68062 800
rect 70030 0 70086 800
rect 72054 0 72110 800
rect 74078 0 74134 800
rect 76102 0 76158 800
rect 78126 0 78182 800
rect 80150 0 80206 800
rect 82174 0 82230 800
rect 84198 0 84254 800
rect 86222 0 86278 800
rect 88246 0 88302 800
rect 90270 0 90326 800
rect 92294 0 92350 800
rect 94318 0 94374 800
rect 96342 0 96398 800
rect 98366 0 98422 800
rect 100390 0 100446 800
rect 102414 0 102470 800
rect 104438 0 104494 800
rect 106462 0 106518 800
rect 108486 0 108542 800
rect 110510 0 110566 800
rect 112534 0 112590 800
rect 114558 0 114614 800
rect 116582 0 116638 800
rect 118606 0 118662 800
rect 120630 0 120686 800
rect 122654 0 122710 800
rect 124678 0 124734 800
rect 126702 0 126758 800
rect 128726 0 128782 800
rect 130750 0 130806 800
rect 132774 0 132830 800
<< obsm2 >>
rect 1216 135456 2354 135674
rect 2522 135456 4010 135674
rect 4178 135456 5666 135674
rect 5834 135456 7322 135674
rect 7490 135456 8978 135674
rect 9146 135456 10634 135674
rect 10802 135456 12290 135674
rect 12458 135456 13946 135674
rect 14114 135456 15602 135674
rect 15770 135456 17258 135674
rect 17426 135456 18914 135674
rect 19082 135456 20570 135674
rect 20738 135456 22226 135674
rect 22394 135456 23882 135674
rect 24050 135456 25538 135674
rect 25706 135456 27194 135674
rect 27362 135456 28850 135674
rect 29018 135456 30506 135674
rect 30674 135456 32162 135674
rect 32330 135456 33818 135674
rect 33986 135456 35474 135674
rect 35642 135456 37130 135674
rect 37298 135456 38786 135674
rect 38954 135456 40442 135674
rect 40610 135456 42098 135674
rect 42266 135456 43754 135674
rect 43922 135456 45410 135674
rect 45578 135456 47066 135674
rect 47234 135456 48722 135674
rect 48890 135456 50378 135674
rect 50546 135456 52034 135674
rect 52202 135456 53690 135674
rect 53858 135456 55346 135674
rect 55514 135456 57002 135674
rect 57170 135456 58658 135674
rect 58826 135456 60314 135674
rect 60482 135456 61970 135674
rect 62138 135456 63626 135674
rect 63794 135456 65282 135674
rect 65450 135456 66938 135674
rect 67106 135456 68594 135674
rect 68762 135456 70250 135674
rect 70418 135456 71906 135674
rect 72074 135456 73562 135674
rect 73730 135456 75218 135674
rect 75386 135456 76874 135674
rect 77042 135456 78530 135674
rect 78698 135456 80186 135674
rect 80354 135456 81842 135674
rect 82010 135456 83498 135674
rect 83666 135456 85154 135674
rect 85322 135456 86810 135674
rect 86978 135456 88466 135674
rect 88634 135456 90122 135674
rect 90290 135456 91778 135674
rect 91946 135456 93434 135674
rect 93602 135456 95090 135674
rect 95258 135456 96746 135674
rect 96914 135456 98402 135674
rect 98570 135456 100058 135674
rect 100226 135456 101714 135674
rect 101882 135456 103370 135674
rect 103538 135456 105026 135674
rect 105194 135456 106682 135674
rect 106850 135456 108338 135674
rect 108506 135456 109994 135674
rect 110162 135456 111650 135674
rect 111818 135456 113306 135674
rect 113474 135456 114962 135674
rect 115130 135456 116618 135674
rect 116786 135456 118274 135674
rect 118442 135456 119930 135674
rect 120098 135456 121586 135674
rect 121754 135456 123242 135674
rect 123410 135456 124898 135674
rect 125066 135456 126554 135674
rect 126722 135456 128210 135674
rect 128378 135456 129866 135674
rect 130034 135456 131522 135674
rect 131690 135456 132816 135674
rect 1216 856 132816 135456
rect 1326 734 3182 856
rect 3350 734 5206 856
rect 5374 734 7230 856
rect 7398 734 9254 856
rect 9422 734 11278 856
rect 11446 734 13302 856
rect 13470 734 15326 856
rect 15494 734 17350 856
rect 17518 734 19374 856
rect 19542 734 21398 856
rect 21566 734 23422 856
rect 23590 734 25446 856
rect 25614 734 27470 856
rect 27638 734 29494 856
rect 29662 734 31518 856
rect 31686 734 33542 856
rect 33710 734 35566 856
rect 35734 734 37590 856
rect 37758 734 39614 856
rect 39782 734 41638 856
rect 41806 734 43662 856
rect 43830 734 45686 856
rect 45854 734 47710 856
rect 47878 734 49734 856
rect 49902 734 51758 856
rect 51926 734 53782 856
rect 53950 734 55806 856
rect 55974 734 57830 856
rect 57998 734 59854 856
rect 60022 734 61878 856
rect 62046 734 63902 856
rect 64070 734 65926 856
rect 66094 734 67950 856
rect 68118 734 69974 856
rect 70142 734 71998 856
rect 72166 734 74022 856
rect 74190 734 76046 856
rect 76214 734 78070 856
rect 78238 734 80094 856
rect 80262 734 82118 856
rect 82286 734 84142 856
rect 84310 734 86166 856
rect 86334 734 88190 856
rect 88358 734 90214 856
rect 90382 734 92238 856
rect 92406 734 94262 856
rect 94430 734 96286 856
rect 96454 734 98310 856
rect 98478 734 100334 856
rect 100502 734 102358 856
rect 102526 734 104382 856
rect 104550 734 106406 856
rect 106574 734 108430 856
rect 108598 734 110454 856
rect 110622 734 112478 856
rect 112646 734 114502 856
rect 114670 734 116526 856
rect 116694 734 118550 856
rect 118718 734 120574 856
rect 120742 734 122598 856
rect 122766 734 124622 856
rect 124790 734 126646 856
rect 126814 734 128670 856
rect 128838 734 130694 856
rect 130862 734 132718 856
<< metal3 >>
rect 133368 102008 134168 102128
rect 133368 34008 134168 34128
<< obsm3 >>
rect 2037 102208 133368 133857
rect 2037 101928 133288 102208
rect 2037 34208 133368 101928
rect 2037 33928 133288 34208
rect 2037 2143 133368 33928
<< metal4 >>
rect 4208 2128 4528 133872
rect 19568 2128 19888 133872
rect 34928 2128 35248 133872
rect 50288 2128 50608 133872
rect 65648 2128 65968 133872
rect 81008 2128 81328 133872
rect 96368 2128 96688 133872
rect 111728 2128 112048 133872
rect 127088 2128 127408 133872
<< obsm4 >>
rect 5947 2483 19488 132701
rect 19968 2483 34848 132701
rect 35328 2483 50208 132701
rect 50688 2483 65568 132701
rect 66048 2483 80928 132701
rect 81408 2483 96288 132701
rect 96768 2483 111648 132701
rect 112128 2483 118069 132701
<< labels >>
rlabel metal2 s 18970 135512 19026 136312 6 becStatus[0]
port 1 nsew signal input
rlabel metal2 s 20626 135512 20682 136312 6 becStatus[1]
port 2 nsew signal input
rlabel metal2 s 22282 135512 22338 136312 6 becStatus[2]
port 3 nsew signal input
rlabel metal2 s 23938 135512 23994 136312 6 becStatus[3]
port 4 nsew signal input
rlabel metal2 s 27250 135512 27306 136312 6 data_in[0]
port 5 nsew signal input
rlabel metal2 s 60370 135512 60426 136312 6 data_in[10]
port 6 nsew signal input
rlabel metal2 s 63682 135512 63738 136312 6 data_in[11]
port 7 nsew signal input
rlabel metal2 s 66994 135512 67050 136312 6 data_in[12]
port 8 nsew signal input
rlabel metal2 s 70306 135512 70362 136312 6 data_in[13]
port 9 nsew signal input
rlabel metal2 s 73618 135512 73674 136312 6 data_in[14]
port 10 nsew signal input
rlabel metal2 s 76930 135512 76986 136312 6 data_in[15]
port 11 nsew signal input
rlabel metal2 s 80242 135512 80298 136312 6 data_in[16]
port 12 nsew signal input
rlabel metal2 s 83554 135512 83610 136312 6 data_in[17]
port 13 nsew signal input
rlabel metal2 s 86866 135512 86922 136312 6 data_in[18]
port 14 nsew signal input
rlabel metal2 s 90178 135512 90234 136312 6 data_in[19]
port 15 nsew signal input
rlabel metal2 s 30562 135512 30618 136312 6 data_in[1]
port 16 nsew signal input
rlabel metal2 s 93490 135512 93546 136312 6 data_in[20]
port 17 nsew signal input
rlabel metal2 s 96802 135512 96858 136312 6 data_in[21]
port 18 nsew signal input
rlabel metal2 s 100114 135512 100170 136312 6 data_in[22]
port 19 nsew signal input
rlabel metal2 s 103426 135512 103482 136312 6 data_in[23]
port 20 nsew signal input
rlabel metal2 s 106738 135512 106794 136312 6 data_in[24]
port 21 nsew signal input
rlabel metal2 s 110050 135512 110106 136312 6 data_in[25]
port 22 nsew signal input
rlabel metal2 s 113362 135512 113418 136312 6 data_in[26]
port 23 nsew signal input
rlabel metal2 s 116674 135512 116730 136312 6 data_in[27]
port 24 nsew signal input
rlabel metal2 s 119986 135512 120042 136312 6 data_in[28]
port 25 nsew signal input
rlabel metal2 s 123298 135512 123354 136312 6 data_in[29]
port 26 nsew signal input
rlabel metal2 s 33874 135512 33930 136312 6 data_in[2]
port 27 nsew signal input
rlabel metal2 s 126610 135512 126666 136312 6 data_in[30]
port 28 nsew signal input
rlabel metal2 s 129922 135512 129978 136312 6 data_in[31]
port 29 nsew signal input
rlabel metal2 s 37186 135512 37242 136312 6 data_in[3]
port 30 nsew signal input
rlabel metal2 s 40498 135512 40554 136312 6 data_in[4]
port 31 nsew signal input
rlabel metal2 s 43810 135512 43866 136312 6 data_in[5]
port 32 nsew signal input
rlabel metal2 s 47122 135512 47178 136312 6 data_in[6]
port 33 nsew signal input
rlabel metal2 s 50434 135512 50490 136312 6 data_in[7]
port 34 nsew signal input
rlabel metal2 s 53746 135512 53802 136312 6 data_in[8]
port 35 nsew signal input
rlabel metal2 s 57058 135512 57114 136312 6 data_in[9]
port 36 nsew signal input
rlabel metal2 s 28906 135512 28962 136312 6 data_out[0]
port 37 nsew signal output
rlabel metal2 s 62026 135512 62082 136312 6 data_out[10]
port 38 nsew signal output
rlabel metal2 s 65338 135512 65394 136312 6 data_out[11]
port 39 nsew signal output
rlabel metal2 s 68650 135512 68706 136312 6 data_out[12]
port 40 nsew signal output
rlabel metal2 s 71962 135512 72018 136312 6 data_out[13]
port 41 nsew signal output
rlabel metal2 s 75274 135512 75330 136312 6 data_out[14]
port 42 nsew signal output
rlabel metal2 s 78586 135512 78642 136312 6 data_out[15]
port 43 nsew signal output
rlabel metal2 s 81898 135512 81954 136312 6 data_out[16]
port 44 nsew signal output
rlabel metal2 s 85210 135512 85266 136312 6 data_out[17]
port 45 nsew signal output
rlabel metal2 s 88522 135512 88578 136312 6 data_out[18]
port 46 nsew signal output
rlabel metal2 s 91834 135512 91890 136312 6 data_out[19]
port 47 nsew signal output
rlabel metal2 s 32218 135512 32274 136312 6 data_out[1]
port 48 nsew signal output
rlabel metal2 s 95146 135512 95202 136312 6 data_out[20]
port 49 nsew signal output
rlabel metal2 s 98458 135512 98514 136312 6 data_out[21]
port 50 nsew signal output
rlabel metal2 s 101770 135512 101826 136312 6 data_out[22]
port 51 nsew signal output
rlabel metal2 s 105082 135512 105138 136312 6 data_out[23]
port 52 nsew signal output
rlabel metal2 s 108394 135512 108450 136312 6 data_out[24]
port 53 nsew signal output
rlabel metal2 s 111706 135512 111762 136312 6 data_out[25]
port 54 nsew signal output
rlabel metal2 s 115018 135512 115074 136312 6 data_out[26]
port 55 nsew signal output
rlabel metal2 s 118330 135512 118386 136312 6 data_out[27]
port 56 nsew signal output
rlabel metal2 s 121642 135512 121698 136312 6 data_out[28]
port 57 nsew signal output
rlabel metal2 s 124954 135512 125010 136312 6 data_out[29]
port 58 nsew signal output
rlabel metal2 s 35530 135512 35586 136312 6 data_out[2]
port 59 nsew signal output
rlabel metal2 s 128266 135512 128322 136312 6 data_out[30]
port 60 nsew signal output
rlabel metal2 s 131578 135512 131634 136312 6 data_out[31]
port 61 nsew signal output
rlabel metal2 s 38842 135512 38898 136312 6 data_out[3]
port 62 nsew signal output
rlabel metal2 s 42154 135512 42210 136312 6 data_out[4]
port 63 nsew signal output
rlabel metal2 s 45466 135512 45522 136312 6 data_out[5]
port 64 nsew signal output
rlabel metal2 s 48778 135512 48834 136312 6 data_out[6]
port 65 nsew signal output
rlabel metal2 s 52090 135512 52146 136312 6 data_out[7]
port 66 nsew signal output
rlabel metal2 s 55402 135512 55458 136312 6 data_out[8]
port 67 nsew signal output
rlabel metal2 s 58714 135512 58770 136312 6 data_out[9]
port 68 nsew signal output
rlabel metal3 s 133368 102008 134168 102128 6 io_oeb
port 69 nsew signal output
rlabel metal3 s 133368 34008 134168 34128 6 io_out
port 70 nsew signal output
rlabel metal2 s 14002 135512 14058 136312 6 ki
port 71 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 la_data_in[0]
port 72 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[10]
port 73 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[11]
port 74 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[12]
port 75 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[13]
port 76 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[14]
port 77 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[15]
port 78 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[16]
port 79 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[17]
port 80 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[18]
port 81 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[19]
port 82 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 la_data_in[1]
port 83 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[20]
port 84 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[21]
port 85 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[22]
port 86 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[23]
port 87 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[24]
port 88 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[25]
port 89 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[26]
port 90 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[27]
port 91 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[28]
port 92 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[29]
port 93 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 la_data_in[2]
port 94 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[30]
port 95 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[31]
port 96 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_data_in[3]
port 97 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 la_data_in[4]
port 98 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_data_in[5]
port 99 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[6]
port 100 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[7]
port 101 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in[8]
port 102 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[9]
port 103 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 la_data_out[0]
port 104 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[10]
port 105 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[11]
port 106 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[12]
port 107 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[13]
port 108 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[14]
port 109 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[15]
port 110 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[16]
port 111 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[17]
port 112 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[18]
port 113 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[19]
port 114 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 la_data_out[1]
port 115 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[20]
port 116 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[21]
port 117 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[22]
port 118 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[23]
port 119 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[24]
port 120 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[25]
port 121 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[26]
port 122 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[27]
port 123 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 la_data_out[28]
port 124 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[29]
port 125 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 la_data_out[2]
port 126 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[30]
port 127 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[31]
port 128 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 la_data_out[3]
port 129 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[4]
port 130 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[5]
port 131 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[6]
port 132 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[7]
port 133 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[8]
port 134 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[9]
port 135 nsew signal output
rlabel metal2 s 12346 135512 12402 136312 6 load_data
port 136 nsew signal output
rlabel metal2 s 2410 135512 2466 136312 6 load_status[0]
port 137 nsew signal output
rlabel metal2 s 4066 135512 4122 136312 6 load_status[1]
port 138 nsew signal output
rlabel metal2 s 5722 135512 5778 136312 6 load_status[2]
port 139 nsew signal output
rlabel metal2 s 7378 135512 7434 136312 6 load_status[3]
port 140 nsew signal output
rlabel metal2 s 9034 135512 9090 136312 6 load_status[4]
port 141 nsew signal output
rlabel metal2 s 10690 135512 10746 136312 6 load_status[5]
port 142 nsew signal output
rlabel metal2 s 15658 135512 15714 136312 6 next_key
port 143 nsew signal input
rlabel metal2 s 17314 135512 17370 136312 6 slv_done
port 144 nsew signal input
rlabel metal2 s 25594 135512 25650 136312 6 slv_enable
port 145 nsew signal output
rlabel metal4 s 4208 2128 4528 133872 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 133872 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 133872 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 133872 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 133872 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 133872 6 vssd1
port 147 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 133872 6 vssd1
port 147 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 133872 6 vssd1
port 147 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 133872 6 vssd1
port 147 nsew ground bidirectional
rlabel metal2 s 1214 0 1270 800 6 wb_clk_i
port 148 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wb_rst_i
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 134168 136312
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 39209060
string GDS_FILE /home/admin/projects/IC5-CASS-2024_2/openlane/lovers_controller/runs/24_11_11_11_05/results/signoff/lovers_controller.magic.gds
string GDS_START 627706
<< end >>

