VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ascon_wrapper
  CLASS BLOCK ;
  FOREIGN ascon_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 449.050 596.000 449.330 600.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 568.520 600.000 569.120 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 470.600 600.000 471.200 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 372.680 600.000 373.280 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 274.760 600.000 275.360 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 176.840 600.000 177.440 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 78.920 600.000 79.520 ;
    END
  END io_in[5]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 596.000 269.930 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 596.000 389.530 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 596.000 150.330 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 596.000 30.730 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 519.560 600.000 520.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 421.640 600.000 422.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 323.720 600.000 324.320 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 225.800 600.000 226.400 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 127.880 600.000 128.480 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 29.960 600.000 30.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 596.000 509.130 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 596.000 329.730 600.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 596.000 210.130 600.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 596.000 90.530 600.000 ;
    END
  END io_out[2]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 596.000 568.930 600.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 594.510 586.215 ;
        RECT 5.330 577.945 594.510 580.775 ;
        RECT 5.330 572.505 594.510 575.335 ;
        RECT 5.330 567.065 594.510 569.895 ;
        RECT 5.330 561.625 594.510 564.455 ;
        RECT 5.330 556.185 594.510 559.015 ;
        RECT 5.330 550.745 594.510 553.575 ;
        RECT 5.330 545.305 594.510 548.135 ;
        RECT 5.330 539.865 594.510 542.695 ;
        RECT 5.330 534.425 594.510 537.255 ;
        RECT 5.330 528.985 594.510 531.815 ;
        RECT 5.330 523.545 594.510 526.375 ;
        RECT 5.330 518.105 594.510 520.935 ;
        RECT 5.330 512.665 594.510 515.495 ;
        RECT 5.330 507.225 594.510 510.055 ;
        RECT 5.330 501.785 594.510 504.615 ;
        RECT 5.330 496.345 594.510 499.175 ;
        RECT 5.330 490.905 594.510 493.735 ;
        RECT 5.330 485.465 594.510 488.295 ;
        RECT 5.330 480.025 594.510 482.855 ;
        RECT 5.330 474.585 594.510 477.415 ;
        RECT 5.330 469.145 594.510 471.975 ;
        RECT 5.330 463.705 594.510 466.535 ;
        RECT 5.330 458.265 594.510 461.095 ;
        RECT 5.330 452.825 594.510 455.655 ;
        RECT 5.330 447.385 594.510 450.215 ;
        RECT 5.330 441.945 594.510 444.775 ;
        RECT 5.330 436.505 594.510 439.335 ;
        RECT 5.330 431.065 594.510 433.895 ;
        RECT 5.330 425.625 594.510 428.455 ;
        RECT 5.330 420.185 594.510 423.015 ;
        RECT 5.330 414.745 594.510 417.575 ;
        RECT 5.330 409.305 594.510 412.135 ;
        RECT 5.330 403.865 594.510 406.695 ;
        RECT 5.330 398.425 594.510 401.255 ;
        RECT 5.330 392.985 594.510 395.815 ;
        RECT 5.330 387.545 594.510 390.375 ;
        RECT 5.330 382.105 594.510 384.935 ;
        RECT 5.330 376.665 594.510 379.495 ;
        RECT 5.330 371.225 594.510 374.055 ;
        RECT 5.330 365.785 594.510 368.615 ;
        RECT 5.330 360.345 594.510 363.175 ;
        RECT 5.330 354.905 594.510 357.735 ;
        RECT 5.330 349.465 594.510 352.295 ;
        RECT 5.330 344.025 594.510 346.855 ;
        RECT 5.330 338.585 594.510 341.415 ;
        RECT 5.330 333.145 594.510 335.975 ;
        RECT 5.330 327.705 594.510 330.535 ;
        RECT 5.330 322.265 594.510 325.095 ;
        RECT 5.330 316.825 594.510 319.655 ;
        RECT 5.330 311.385 594.510 314.215 ;
        RECT 5.330 305.945 594.510 308.775 ;
        RECT 5.330 300.505 594.510 303.335 ;
        RECT 5.330 295.065 594.510 297.895 ;
        RECT 5.330 289.625 594.510 292.455 ;
        RECT 5.330 284.185 594.510 287.015 ;
        RECT 5.330 278.745 594.510 281.575 ;
        RECT 5.330 273.305 594.510 276.135 ;
        RECT 5.330 267.865 594.510 270.695 ;
        RECT 5.330 262.425 594.510 265.255 ;
        RECT 5.330 256.985 594.510 259.815 ;
        RECT 5.330 251.545 594.510 254.375 ;
        RECT 5.330 246.105 594.510 248.935 ;
        RECT 5.330 240.665 594.510 243.495 ;
        RECT 5.330 235.225 594.510 238.055 ;
        RECT 5.330 229.785 594.510 232.615 ;
        RECT 5.330 224.345 594.510 227.175 ;
        RECT 5.330 218.905 594.510 221.735 ;
        RECT 5.330 213.465 594.510 216.295 ;
        RECT 5.330 208.025 594.510 210.855 ;
        RECT 5.330 202.585 594.510 205.415 ;
        RECT 5.330 197.145 594.510 199.975 ;
        RECT 5.330 191.705 594.510 194.535 ;
        RECT 5.330 186.265 594.510 189.095 ;
        RECT 5.330 180.825 594.510 183.655 ;
        RECT 5.330 175.385 594.510 178.215 ;
        RECT 5.330 169.945 594.510 172.775 ;
        RECT 5.330 164.505 594.510 167.335 ;
        RECT 5.330 159.065 594.510 161.895 ;
        RECT 5.330 153.625 594.510 156.455 ;
        RECT 5.330 148.185 594.510 151.015 ;
        RECT 5.330 142.745 594.510 145.575 ;
        RECT 5.330 137.305 594.510 140.135 ;
        RECT 5.330 131.865 594.510 134.695 ;
        RECT 5.330 126.425 594.510 129.255 ;
        RECT 5.330 120.985 594.510 123.815 ;
        RECT 5.330 115.545 594.510 118.375 ;
        RECT 5.330 110.105 594.510 112.935 ;
        RECT 5.330 104.665 594.510 107.495 ;
        RECT 5.330 99.225 594.510 102.055 ;
        RECT 5.330 93.785 594.510 96.615 ;
        RECT 5.330 88.345 594.510 91.175 ;
        RECT 5.330 82.905 594.510 85.735 ;
        RECT 5.330 77.465 594.510 80.295 ;
        RECT 5.330 72.025 594.510 74.855 ;
        RECT 5.330 66.585 594.510 69.415 ;
        RECT 5.330 61.145 594.510 63.975 ;
        RECT 5.330 55.705 594.510 58.535 ;
        RECT 5.330 50.265 594.510 53.095 ;
        RECT 5.330 44.825 594.510 47.655 ;
        RECT 5.330 39.385 594.510 42.215 ;
        RECT 5.330 33.945 594.510 36.775 ;
        RECT 5.330 28.505 594.510 31.335 ;
        RECT 5.330 23.065 594.510 25.895 ;
        RECT 5.330 17.625 594.510 20.455 ;
        RECT 5.330 12.185 594.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 594.620 587.760 ;
      LAYER met2 ;
        RECT 7.000 595.720 30.170 596.770 ;
        RECT 31.010 595.720 89.970 596.770 ;
        RECT 90.810 595.720 149.770 596.770 ;
        RECT 150.610 595.720 209.570 596.770 ;
        RECT 210.410 595.720 269.370 596.770 ;
        RECT 270.210 595.720 329.170 596.770 ;
        RECT 330.010 595.720 388.970 596.770 ;
        RECT 389.810 595.720 448.770 596.770 ;
        RECT 449.610 595.720 508.570 596.770 ;
        RECT 509.410 595.720 568.370 596.770 ;
        RECT 569.210 595.720 594.230 596.770 ;
        RECT 7.000 10.695 594.230 595.720 ;
      LAYER met3 ;
        RECT 10.645 569.520 596.000 587.685 ;
        RECT 10.645 568.120 595.600 569.520 ;
        RECT 10.645 520.560 596.000 568.120 ;
        RECT 10.645 519.160 595.600 520.560 ;
        RECT 10.645 471.600 596.000 519.160 ;
        RECT 10.645 470.200 595.600 471.600 ;
        RECT 10.645 422.640 596.000 470.200 ;
        RECT 10.645 421.240 595.600 422.640 ;
        RECT 10.645 373.680 596.000 421.240 ;
        RECT 10.645 372.280 595.600 373.680 ;
        RECT 10.645 324.720 596.000 372.280 ;
        RECT 10.645 323.320 595.600 324.720 ;
        RECT 10.645 275.760 596.000 323.320 ;
        RECT 10.645 274.360 595.600 275.760 ;
        RECT 10.645 226.800 596.000 274.360 ;
        RECT 10.645 225.400 595.600 226.800 ;
        RECT 10.645 177.840 596.000 225.400 ;
        RECT 10.645 176.440 595.600 177.840 ;
        RECT 10.645 128.880 596.000 176.440 ;
        RECT 10.645 127.480 595.600 128.880 ;
        RECT 10.645 79.920 596.000 127.480 ;
        RECT 10.645 78.520 595.600 79.920 ;
        RECT 10.645 30.960 596.000 78.520 ;
        RECT 10.645 29.560 595.600 30.960 ;
        RECT 10.645 10.715 596.000 29.560 ;
      LAYER met4 ;
        RECT 11.335 27.375 20.640 573.065 ;
        RECT 23.040 27.375 97.440 573.065 ;
        RECT 99.840 27.375 174.240 573.065 ;
        RECT 176.640 27.375 251.040 573.065 ;
        RECT 253.440 27.375 327.840 573.065 ;
        RECT 330.240 27.375 404.640 573.065 ;
        RECT 407.040 27.375 481.440 573.065 ;
        RECT 483.840 27.375 558.240 573.065 ;
        RECT 560.640 27.375 575.625 573.065 ;
  END
END ascon_wrapper
END LIBRARY

