VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lovers_controller
  CLASS BLOCK ;
  FOREIGN lovers_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 670.840 BY 681.560 ;
  PIN becStatus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 677.560 95.130 681.560 ;
    END
  END becStatus[0]
  PIN becStatus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 677.560 103.410 681.560 ;
    END
  END becStatus[1]
  PIN becStatus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 677.560 111.690 681.560 ;
    END
  END becStatus[2]
  PIN becStatus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 677.560 119.970 681.560 ;
    END
  END becStatus[3]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 136.250 677.560 136.530 681.560 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 301.850 677.560 302.130 681.560 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 677.560 318.690 681.560 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 677.560 335.250 681.560 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 351.530 677.560 351.810 681.560 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 677.560 368.370 681.560 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 384.650 677.560 384.930 681.560 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 401.210 677.560 401.490 681.560 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 417.770 677.560 418.050 681.560 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 434.330 677.560 434.610 681.560 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 450.890 677.560 451.170 681.560 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 152.810 677.560 153.090 681.560 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 467.450 677.560 467.730 681.560 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 677.560 484.290 681.560 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 500.570 677.560 500.850 681.560 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 517.130 677.560 517.410 681.560 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 533.690 677.560 533.970 681.560 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 550.250 677.560 550.530 681.560 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 566.810 677.560 567.090 681.560 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 583.370 677.560 583.650 681.560 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 599.930 677.560 600.210 681.560 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 616.490 677.560 616.770 681.560 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 677.560 169.650 681.560 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 633.050 677.560 633.330 681.560 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 649.610 677.560 649.890 681.560 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 185.930 677.560 186.210 681.560 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 202.490 677.560 202.770 681.560 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 677.560 219.330 681.560 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.610 677.560 235.890 681.560 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 252.170 677.560 252.450 681.560 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 677.560 269.010 681.560 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 285.290 677.560 285.570 681.560 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 677.560 144.810 681.560 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 677.560 310.410 681.560 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 326.690 677.560 326.970 681.560 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 677.560 343.530 681.560 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 359.810 677.560 360.090 681.560 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 376.370 677.560 376.650 681.560 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 677.560 393.210 681.560 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 677.560 409.770 681.560 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 426.050 677.560 426.330 681.560 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 442.610 677.560 442.890 681.560 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 459.170 677.560 459.450 681.560 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 677.560 161.370 681.560 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 475.730 677.560 476.010 681.560 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 492.290 677.560 492.570 681.560 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 508.850 677.560 509.130 681.560 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 525.410 677.560 525.690 681.560 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 541.970 677.560 542.250 681.560 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 558.530 677.560 558.810 681.560 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 677.560 575.370 681.560 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 591.650 677.560 591.930 681.560 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 608.210 677.560 608.490 681.560 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 624.770 677.560 625.050 681.560 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 677.560 177.930 681.560 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 641.330 677.560 641.610 681.560 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 657.890 677.560 658.170 681.560 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 677.560 194.490 681.560 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 677.560 211.050 681.560 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 227.330 677.560 227.610 681.560 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 677.560 244.170 681.560 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 677.560 260.730 681.560 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 677.560 277.290 681.560 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 677.560 293.850 681.560 ;
    END
  END data_out[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 666.840 510.040 670.840 510.640 ;
    END
  END io_oeb
  PIN io_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 666.840 170.040 670.840 170.640 ;
    END
  END io_out
  PIN ki
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 677.560 70.290 681.560 ;
    END
  END ki
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la_data_out[9]
  PIN load_data
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 677.560 62.010 681.560 ;
    END
  END load_data
  PIN load_status[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 12.050 677.560 12.330 681.560 ;
    END
  END load_status[0]
  PIN load_status[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 677.560 20.610 681.560 ;
    END
  END load_status[1]
  PIN load_status[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 677.560 28.890 681.560 ;
    END
  END load_status[2]
  PIN load_status[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 677.560 37.170 681.560 ;
    END
  END load_status[3]
  PIN load_status[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 677.560 45.450 681.560 ;
    END
  END load_status[4]
  PIN load_status[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 53.450 677.560 53.730 681.560 ;
    END
  END load_status[5]
  PIN next_key
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 677.560 78.570 681.560 ;
    END
  END next_key
  PIN slv_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 86.570 677.560 86.850 681.560 ;
    END
  END slv_done
  PIN slv_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 677.560 128.250 681.560 ;
    END
  END slv_enable
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 669.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 669.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 669.360 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 664.985 665.350 667.815 ;
        RECT 5.330 659.545 665.350 662.375 ;
        RECT 5.330 654.105 665.350 656.935 ;
        RECT 5.330 648.665 665.350 651.495 ;
        RECT 5.330 643.225 665.350 646.055 ;
        RECT 5.330 637.785 665.350 640.615 ;
        RECT 5.330 632.345 665.350 635.175 ;
        RECT 5.330 626.905 665.350 629.735 ;
        RECT 5.330 621.465 665.350 624.295 ;
        RECT 5.330 616.025 665.350 618.855 ;
        RECT 5.330 610.585 665.350 613.415 ;
        RECT 5.330 605.145 665.350 607.975 ;
        RECT 5.330 599.705 665.350 602.535 ;
        RECT 5.330 594.265 665.350 597.095 ;
        RECT 5.330 588.825 665.350 591.655 ;
        RECT 5.330 583.385 665.350 586.215 ;
        RECT 5.330 577.945 665.350 580.775 ;
        RECT 5.330 572.505 665.350 575.335 ;
        RECT 5.330 567.065 665.350 569.895 ;
        RECT 5.330 561.625 665.350 564.455 ;
        RECT 5.330 556.185 665.350 559.015 ;
        RECT 5.330 550.745 665.350 553.575 ;
        RECT 5.330 545.305 665.350 548.135 ;
        RECT 5.330 539.865 665.350 542.695 ;
        RECT 5.330 534.425 665.350 537.255 ;
        RECT 5.330 528.985 665.350 531.815 ;
        RECT 5.330 523.545 665.350 526.375 ;
        RECT 5.330 518.105 665.350 520.935 ;
        RECT 5.330 512.665 665.350 515.495 ;
        RECT 5.330 507.225 665.350 510.055 ;
        RECT 5.330 501.785 665.350 504.615 ;
        RECT 5.330 496.345 665.350 499.175 ;
        RECT 5.330 490.905 665.350 493.735 ;
        RECT 5.330 485.465 665.350 488.295 ;
        RECT 5.330 480.025 665.350 482.855 ;
        RECT 5.330 474.585 665.350 477.415 ;
        RECT 5.330 469.145 665.350 471.975 ;
        RECT 5.330 463.705 665.350 466.535 ;
        RECT 5.330 458.265 665.350 461.095 ;
        RECT 5.330 452.825 665.350 455.655 ;
        RECT 5.330 447.385 665.350 450.215 ;
        RECT 5.330 441.945 665.350 444.775 ;
        RECT 5.330 436.505 665.350 439.335 ;
        RECT 5.330 431.065 665.350 433.895 ;
        RECT 5.330 425.625 665.350 428.455 ;
        RECT 5.330 420.185 665.350 423.015 ;
        RECT 5.330 414.745 665.350 417.575 ;
        RECT 5.330 409.305 665.350 412.135 ;
        RECT 5.330 403.865 665.350 406.695 ;
        RECT 5.330 398.425 665.350 401.255 ;
        RECT 5.330 392.985 665.350 395.815 ;
        RECT 5.330 387.545 665.350 390.375 ;
        RECT 5.330 382.105 665.350 384.935 ;
        RECT 5.330 376.665 665.350 379.495 ;
        RECT 5.330 371.225 665.350 374.055 ;
        RECT 5.330 365.785 665.350 368.615 ;
        RECT 5.330 360.345 665.350 363.175 ;
        RECT 5.330 354.905 665.350 357.735 ;
        RECT 5.330 349.465 665.350 352.295 ;
        RECT 5.330 344.025 665.350 346.855 ;
        RECT 5.330 338.585 665.350 341.415 ;
        RECT 5.330 333.145 665.350 335.975 ;
        RECT 5.330 327.705 665.350 330.535 ;
        RECT 5.330 322.265 665.350 325.095 ;
        RECT 5.330 316.825 665.350 319.655 ;
        RECT 5.330 311.385 665.350 314.215 ;
        RECT 5.330 305.945 665.350 308.775 ;
        RECT 5.330 300.505 665.350 303.335 ;
        RECT 5.330 295.065 665.350 297.895 ;
        RECT 5.330 289.625 665.350 292.455 ;
        RECT 5.330 284.185 665.350 287.015 ;
        RECT 5.330 278.745 665.350 281.575 ;
        RECT 5.330 273.305 665.350 276.135 ;
        RECT 5.330 267.865 665.350 270.695 ;
        RECT 5.330 262.425 665.350 265.255 ;
        RECT 5.330 256.985 665.350 259.815 ;
        RECT 5.330 251.545 665.350 254.375 ;
        RECT 5.330 246.105 665.350 248.935 ;
        RECT 5.330 240.665 665.350 243.495 ;
        RECT 5.330 235.225 665.350 238.055 ;
        RECT 5.330 229.785 665.350 232.615 ;
        RECT 5.330 224.345 665.350 227.175 ;
        RECT 5.330 218.905 665.350 221.735 ;
        RECT 5.330 213.465 665.350 216.295 ;
        RECT 5.330 208.025 665.350 210.855 ;
        RECT 5.330 202.585 665.350 205.415 ;
        RECT 5.330 197.145 665.350 199.975 ;
        RECT 5.330 191.705 665.350 194.535 ;
        RECT 5.330 186.265 665.350 189.095 ;
        RECT 5.330 180.825 665.350 183.655 ;
        RECT 5.330 175.385 665.350 178.215 ;
        RECT 5.330 169.945 665.350 172.775 ;
        RECT 5.330 164.505 665.350 167.335 ;
        RECT 5.330 159.065 665.350 161.895 ;
        RECT 5.330 153.625 665.350 156.455 ;
        RECT 5.330 148.185 665.350 151.015 ;
        RECT 5.330 142.745 665.350 145.575 ;
        RECT 5.330 137.305 665.350 140.135 ;
        RECT 5.330 131.865 665.350 134.695 ;
        RECT 5.330 126.425 665.350 129.255 ;
        RECT 5.330 120.985 665.350 123.815 ;
        RECT 5.330 115.545 665.350 118.375 ;
        RECT 5.330 110.105 665.350 112.935 ;
        RECT 5.330 104.665 665.350 107.495 ;
        RECT 5.330 99.225 665.350 102.055 ;
        RECT 5.330 93.785 665.350 96.615 ;
        RECT 5.330 88.345 665.350 91.175 ;
        RECT 5.330 82.905 665.350 85.735 ;
        RECT 5.330 77.465 665.350 80.295 ;
        RECT 5.330 72.025 665.350 74.855 ;
        RECT 5.330 66.585 665.350 69.415 ;
        RECT 5.330 61.145 665.350 63.975 ;
        RECT 5.330 55.705 665.350 58.535 ;
        RECT 5.330 50.265 665.350 53.095 ;
        RECT 5.330 44.825 665.350 47.655 ;
        RECT 5.330 39.385 665.350 42.215 ;
        RECT 5.330 33.945 665.350 36.775 ;
        RECT 5.330 28.505 665.350 31.335 ;
        RECT 5.330 23.065 665.350 25.895 ;
        RECT 5.330 17.625 665.350 20.455 ;
        RECT 5.330 12.185 665.350 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 665.160 669.205 ;
      LAYER met1 ;
        RECT 5.520 8.880 665.160 669.360 ;
      LAYER met2 ;
        RECT 6.080 677.280 11.770 678.370 ;
        RECT 12.610 677.280 20.050 678.370 ;
        RECT 20.890 677.280 28.330 678.370 ;
        RECT 29.170 677.280 36.610 678.370 ;
        RECT 37.450 677.280 44.890 678.370 ;
        RECT 45.730 677.280 53.170 678.370 ;
        RECT 54.010 677.280 61.450 678.370 ;
        RECT 62.290 677.280 69.730 678.370 ;
        RECT 70.570 677.280 78.010 678.370 ;
        RECT 78.850 677.280 86.290 678.370 ;
        RECT 87.130 677.280 94.570 678.370 ;
        RECT 95.410 677.280 102.850 678.370 ;
        RECT 103.690 677.280 111.130 678.370 ;
        RECT 111.970 677.280 119.410 678.370 ;
        RECT 120.250 677.280 127.690 678.370 ;
        RECT 128.530 677.280 135.970 678.370 ;
        RECT 136.810 677.280 144.250 678.370 ;
        RECT 145.090 677.280 152.530 678.370 ;
        RECT 153.370 677.280 160.810 678.370 ;
        RECT 161.650 677.280 169.090 678.370 ;
        RECT 169.930 677.280 177.370 678.370 ;
        RECT 178.210 677.280 185.650 678.370 ;
        RECT 186.490 677.280 193.930 678.370 ;
        RECT 194.770 677.280 202.210 678.370 ;
        RECT 203.050 677.280 210.490 678.370 ;
        RECT 211.330 677.280 218.770 678.370 ;
        RECT 219.610 677.280 227.050 678.370 ;
        RECT 227.890 677.280 235.330 678.370 ;
        RECT 236.170 677.280 243.610 678.370 ;
        RECT 244.450 677.280 251.890 678.370 ;
        RECT 252.730 677.280 260.170 678.370 ;
        RECT 261.010 677.280 268.450 678.370 ;
        RECT 269.290 677.280 276.730 678.370 ;
        RECT 277.570 677.280 285.010 678.370 ;
        RECT 285.850 677.280 293.290 678.370 ;
        RECT 294.130 677.280 301.570 678.370 ;
        RECT 302.410 677.280 309.850 678.370 ;
        RECT 310.690 677.280 318.130 678.370 ;
        RECT 318.970 677.280 326.410 678.370 ;
        RECT 327.250 677.280 334.690 678.370 ;
        RECT 335.530 677.280 342.970 678.370 ;
        RECT 343.810 677.280 351.250 678.370 ;
        RECT 352.090 677.280 359.530 678.370 ;
        RECT 360.370 677.280 367.810 678.370 ;
        RECT 368.650 677.280 376.090 678.370 ;
        RECT 376.930 677.280 384.370 678.370 ;
        RECT 385.210 677.280 392.650 678.370 ;
        RECT 393.490 677.280 400.930 678.370 ;
        RECT 401.770 677.280 409.210 678.370 ;
        RECT 410.050 677.280 417.490 678.370 ;
        RECT 418.330 677.280 425.770 678.370 ;
        RECT 426.610 677.280 434.050 678.370 ;
        RECT 434.890 677.280 442.330 678.370 ;
        RECT 443.170 677.280 450.610 678.370 ;
        RECT 451.450 677.280 458.890 678.370 ;
        RECT 459.730 677.280 467.170 678.370 ;
        RECT 468.010 677.280 475.450 678.370 ;
        RECT 476.290 677.280 483.730 678.370 ;
        RECT 484.570 677.280 492.010 678.370 ;
        RECT 492.850 677.280 500.290 678.370 ;
        RECT 501.130 677.280 508.570 678.370 ;
        RECT 509.410 677.280 516.850 678.370 ;
        RECT 517.690 677.280 525.130 678.370 ;
        RECT 525.970 677.280 533.410 678.370 ;
        RECT 534.250 677.280 541.690 678.370 ;
        RECT 542.530 677.280 549.970 678.370 ;
        RECT 550.810 677.280 558.250 678.370 ;
        RECT 559.090 677.280 566.530 678.370 ;
        RECT 567.370 677.280 574.810 678.370 ;
        RECT 575.650 677.280 583.090 678.370 ;
        RECT 583.930 677.280 591.370 678.370 ;
        RECT 592.210 677.280 599.650 678.370 ;
        RECT 600.490 677.280 607.930 678.370 ;
        RECT 608.770 677.280 616.210 678.370 ;
        RECT 617.050 677.280 624.490 678.370 ;
        RECT 625.330 677.280 632.770 678.370 ;
        RECT 633.610 677.280 641.050 678.370 ;
        RECT 641.890 677.280 649.330 678.370 ;
        RECT 650.170 677.280 657.610 678.370 ;
        RECT 658.450 677.280 664.080 678.370 ;
        RECT 6.080 4.280 664.080 677.280 ;
        RECT 6.630 3.670 15.910 4.280 ;
        RECT 16.750 3.670 26.030 4.280 ;
        RECT 26.870 3.670 36.150 4.280 ;
        RECT 36.990 3.670 46.270 4.280 ;
        RECT 47.110 3.670 56.390 4.280 ;
        RECT 57.230 3.670 66.510 4.280 ;
        RECT 67.350 3.670 76.630 4.280 ;
        RECT 77.470 3.670 86.750 4.280 ;
        RECT 87.590 3.670 96.870 4.280 ;
        RECT 97.710 3.670 106.990 4.280 ;
        RECT 107.830 3.670 117.110 4.280 ;
        RECT 117.950 3.670 127.230 4.280 ;
        RECT 128.070 3.670 137.350 4.280 ;
        RECT 138.190 3.670 147.470 4.280 ;
        RECT 148.310 3.670 157.590 4.280 ;
        RECT 158.430 3.670 167.710 4.280 ;
        RECT 168.550 3.670 177.830 4.280 ;
        RECT 178.670 3.670 187.950 4.280 ;
        RECT 188.790 3.670 198.070 4.280 ;
        RECT 198.910 3.670 208.190 4.280 ;
        RECT 209.030 3.670 218.310 4.280 ;
        RECT 219.150 3.670 228.430 4.280 ;
        RECT 229.270 3.670 238.550 4.280 ;
        RECT 239.390 3.670 248.670 4.280 ;
        RECT 249.510 3.670 258.790 4.280 ;
        RECT 259.630 3.670 268.910 4.280 ;
        RECT 269.750 3.670 279.030 4.280 ;
        RECT 279.870 3.670 289.150 4.280 ;
        RECT 289.990 3.670 299.270 4.280 ;
        RECT 300.110 3.670 309.390 4.280 ;
        RECT 310.230 3.670 319.510 4.280 ;
        RECT 320.350 3.670 329.630 4.280 ;
        RECT 330.470 3.670 339.750 4.280 ;
        RECT 340.590 3.670 349.870 4.280 ;
        RECT 350.710 3.670 359.990 4.280 ;
        RECT 360.830 3.670 370.110 4.280 ;
        RECT 370.950 3.670 380.230 4.280 ;
        RECT 381.070 3.670 390.350 4.280 ;
        RECT 391.190 3.670 400.470 4.280 ;
        RECT 401.310 3.670 410.590 4.280 ;
        RECT 411.430 3.670 420.710 4.280 ;
        RECT 421.550 3.670 430.830 4.280 ;
        RECT 431.670 3.670 440.950 4.280 ;
        RECT 441.790 3.670 451.070 4.280 ;
        RECT 451.910 3.670 461.190 4.280 ;
        RECT 462.030 3.670 471.310 4.280 ;
        RECT 472.150 3.670 481.430 4.280 ;
        RECT 482.270 3.670 491.550 4.280 ;
        RECT 492.390 3.670 501.670 4.280 ;
        RECT 502.510 3.670 511.790 4.280 ;
        RECT 512.630 3.670 521.910 4.280 ;
        RECT 522.750 3.670 532.030 4.280 ;
        RECT 532.870 3.670 542.150 4.280 ;
        RECT 542.990 3.670 552.270 4.280 ;
        RECT 553.110 3.670 562.390 4.280 ;
        RECT 563.230 3.670 572.510 4.280 ;
        RECT 573.350 3.670 582.630 4.280 ;
        RECT 583.470 3.670 592.750 4.280 ;
        RECT 593.590 3.670 602.870 4.280 ;
        RECT 603.710 3.670 612.990 4.280 ;
        RECT 613.830 3.670 623.110 4.280 ;
        RECT 623.950 3.670 633.230 4.280 ;
        RECT 634.070 3.670 643.350 4.280 ;
        RECT 644.190 3.670 653.470 4.280 ;
        RECT 654.310 3.670 663.590 4.280 ;
      LAYER met3 ;
        RECT 10.185 511.040 666.840 669.285 ;
        RECT 10.185 509.640 666.440 511.040 ;
        RECT 10.185 171.040 666.840 509.640 ;
        RECT 10.185 169.640 666.440 171.040 ;
        RECT 10.185 10.715 666.840 169.640 ;
      LAYER met4 ;
        RECT 29.735 12.415 97.440 663.505 ;
        RECT 99.840 12.415 174.240 663.505 ;
        RECT 176.640 12.415 251.040 663.505 ;
        RECT 253.440 12.415 327.840 663.505 ;
        RECT 330.240 12.415 404.640 663.505 ;
        RECT 407.040 12.415 481.440 663.505 ;
        RECT 483.840 12.415 558.240 663.505 ;
        RECT 560.640 12.415 590.345 663.505 ;
  END
END lovers_controller
END LIBRARY

