magic
tech sky130A
magscale 1 2
timestamp 1730980974
<< nwell >>
rect 1066 97093 98846 97414
rect 1066 96005 98846 96571
rect 1066 94917 98846 95483
rect 1066 93829 98846 94395
rect 1066 92741 98846 93307
rect 1066 91653 98846 92219
rect 1066 90565 98846 91131
rect 1066 89477 98846 90043
rect 1066 88389 98846 88955
rect 1066 87301 98846 87867
rect 1066 86213 98846 86779
rect 1066 85125 98846 85691
rect 1066 84037 98846 84603
rect 1066 82949 98846 83515
rect 1066 81861 98846 82427
rect 1066 80773 98846 81339
rect 1066 79685 98846 80251
rect 1066 78597 98846 79163
rect 1066 77509 98846 78075
rect 1066 76421 98846 76987
rect 1066 75333 98846 75899
rect 1066 74245 98846 74811
rect 1066 73157 98846 73723
rect 1066 72069 98846 72635
rect 1066 70981 98846 71547
rect 1066 69893 98846 70459
rect 1066 68805 98846 69371
rect 1066 67717 98846 68283
rect 1066 66629 98846 67195
rect 1066 65541 98846 66107
rect 1066 64453 98846 65019
rect 1066 63365 98846 63931
rect 1066 62277 98846 62843
rect 1066 61189 98846 61755
rect 1066 60101 98846 60667
rect 1066 59013 98846 59579
rect 1066 57925 98846 58491
rect 1066 56837 98846 57403
rect 1066 55749 98846 56315
rect 1066 54661 98846 55227
rect 1066 53573 98846 54139
rect 1066 52485 98846 53051
rect 1066 51397 98846 51963
rect 1066 50309 98846 50875
rect 1066 49221 98846 49787
rect 1066 48133 98846 48699
rect 1066 47045 98846 47611
rect 1066 45957 98846 46523
rect 1066 44869 98846 45435
rect 1066 43781 98846 44347
rect 1066 42693 98846 43259
rect 1066 41605 98846 42171
rect 1066 40517 98846 41083
rect 1066 39429 98846 39995
rect 1066 38341 98846 38907
rect 1066 37253 98846 37819
rect 1066 36165 98846 36731
rect 1066 35077 98846 35643
rect 1066 33989 98846 34555
rect 1066 32901 98846 33467
rect 1066 31813 98846 32379
rect 1066 30725 98846 31291
rect 1066 29637 98846 30203
rect 1066 28549 98846 29115
rect 1066 27461 98846 28027
rect 1066 26373 98846 26939
rect 1066 25285 98846 25851
rect 1066 24197 98846 24763
rect 1066 23109 98846 23675
rect 1066 22021 98846 22587
rect 1066 20933 98846 21499
rect 1066 19845 98846 20411
rect 1066 18757 98846 19323
rect 1066 17669 98846 18235
rect 1066 16581 98846 17147
rect 1066 15493 98846 16059
rect 1066 14405 98846 14971
rect 1066 13317 98846 13883
rect 1066 12229 98846 12795
rect 1066 11141 98846 11707
rect 1066 10053 98846 10619
rect 1066 8965 98846 9531
rect 1066 7877 98846 8443
rect 1066 6789 98846 7355
rect 1066 5701 98846 6267
rect 1066 4613 98846 5179
rect 1066 3525 98846 4091
rect 1066 2437 98846 3003
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< metal2 >>
rect 1490 0 1546 800
rect 4342 0 4398 800
rect 7194 0 7250 800
rect 10046 0 10102 800
rect 12898 0 12954 800
rect 15750 0 15806 800
rect 18602 0 18658 800
rect 21454 0 21510 800
rect 24306 0 24362 800
rect 27158 0 27214 800
rect 30010 0 30066 800
rect 32862 0 32918 800
rect 35714 0 35770 800
rect 38566 0 38622 800
rect 41418 0 41474 800
rect 44270 0 44326 800
rect 47122 0 47178 800
rect 49974 0 50030 800
rect 52826 0 52882 800
rect 55678 0 55734 800
rect 58530 0 58586 800
rect 61382 0 61438 800
rect 64234 0 64290 800
rect 67086 0 67142 800
rect 69938 0 69994 800
rect 72790 0 72846 800
rect 75642 0 75698 800
rect 78494 0 78550 800
rect 81346 0 81402 800
rect 84198 0 84254 800
rect 87050 0 87106 800
rect 89902 0 89958 800
rect 92754 0 92810 800
rect 95606 0 95662 800
rect 98458 0 98514 800
<< obsm2 >>
rect 1492 856 98500 97413
rect 1602 734 4286 856
rect 4454 734 7138 856
rect 7306 734 9990 856
rect 10158 734 12842 856
rect 13010 734 15694 856
rect 15862 734 18546 856
rect 18714 734 21398 856
rect 21566 734 24250 856
rect 24418 734 27102 856
rect 27270 734 29954 856
rect 30122 734 32806 856
rect 32974 734 35658 856
rect 35826 734 38510 856
rect 38678 734 41362 856
rect 41530 734 44214 856
rect 44382 734 47066 856
rect 47234 734 49918 856
rect 50086 734 52770 856
rect 52938 734 55622 856
rect 55790 734 58474 856
rect 58642 734 61326 856
rect 61494 734 64178 856
rect 64346 734 67030 856
rect 67198 734 69882 856
rect 70050 734 72734 856
rect 72902 734 75586 856
rect 75754 734 78438 856
rect 78606 734 81290 856
rect 81458 734 84142 856
rect 84310 734 86994 856
rect 87162 734 89846 856
rect 90014 734 92698 856
rect 92866 734 95550 856
rect 95718 734 98402 856
<< obsm3 >>
rect 4210 2143 96686 97409
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal2 s 10046 0 10102 800 6 a[0]
port 1 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 a[1]
port 2 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 a[2]
port 3 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 a[3]
port 4 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 a[4]
port 5 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 a[5]
port 6 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 a[6]
port 7 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 a[7]
port 8 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 b[0]
port 9 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 b[1]
port 10 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 b[2]
port 11 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 b[3]
port 12 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 b[4]
port 13 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 b[5]
port 14 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 b[6]
port 15 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 b[7]
port 16 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 clk
port 17 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 control
port 18 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 p[0]
port 19 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 p[10]
port 20 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 p[11]
port 21 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 p[12]
port 22 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 p[13]
port 23 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 p[14]
port 24 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 p[15]
port 25 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 p[1]
port 26 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 p[2]
port 27 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 p[3]
port 28 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 p[4]
port 29 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 p[5]
port 30 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 p[6]
port 31 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 p[7]
port 32 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 p[8]
port 33 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 p[9]
port 34 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 rst
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4438474
string GDS_FILE /home/admin/projects/IC5-CASS-2024/openlane/vmsu_8bit/runs/24_11_07_18_57/results/signoff/vmsu_8bit_top.magic.gds
string GDS_START 333016
<< end >>

