VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bec
  CLASS BLOCK ;
  FOREIGN bec ;
  ORIGIN 0.000 0.000 ;
  SIZE 935.205 BY 945.925 ;
  PIN becStatus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END becStatus[0]
  PIN becStatus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END becStatus[1]
  PIN becStatus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END becStatus[2]
  PIN becStatus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END becStatus[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 869.950 0.000 870.230 4.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 4.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END data_out[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END enable
  PIN ki
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END ki
  PIN load_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END load_data
  PIN load_status[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END load_status[0]
  PIN load_status[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END load_status[1]
  PIN load_status[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END load_status[2]
  PIN load_status[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END load_status[3]
  PIN load_status[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END load_status[4]
  PIN load_status[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END load_status[5]
  PIN next_key
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END next_key
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END rst
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 933.200 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 933.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 933.200 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 5.330 931.545 929.850 933.150 ;
        RECT 5.330 926.105 929.850 928.935 ;
        RECT 5.330 920.665 929.850 923.495 ;
        RECT 5.330 915.225 929.850 918.055 ;
        RECT 5.330 909.785 929.850 912.615 ;
        RECT 5.330 904.345 929.850 907.175 ;
        RECT 5.330 898.905 929.850 901.735 ;
        RECT 5.330 893.465 929.850 896.295 ;
        RECT 5.330 888.025 929.850 890.855 ;
        RECT 5.330 882.585 929.850 885.415 ;
        RECT 5.330 877.145 929.850 879.975 ;
        RECT 5.330 871.705 929.850 874.535 ;
        RECT 5.330 866.265 929.850 869.095 ;
        RECT 5.330 860.825 929.850 863.655 ;
        RECT 5.330 855.385 929.850 858.215 ;
        RECT 5.330 849.945 929.850 852.775 ;
        RECT 5.330 844.505 929.850 847.335 ;
        RECT 5.330 839.065 929.850 841.895 ;
        RECT 5.330 833.625 929.850 836.455 ;
        RECT 5.330 828.185 929.850 831.015 ;
        RECT 5.330 822.745 929.850 825.575 ;
        RECT 5.330 817.305 929.850 820.135 ;
        RECT 5.330 811.865 929.850 814.695 ;
        RECT 5.330 806.425 929.850 809.255 ;
        RECT 5.330 800.985 929.850 803.815 ;
        RECT 5.330 795.545 929.850 798.375 ;
        RECT 5.330 790.105 929.850 792.935 ;
        RECT 5.330 784.665 929.850 787.495 ;
        RECT 5.330 779.225 929.850 782.055 ;
        RECT 5.330 773.785 929.850 776.615 ;
        RECT 5.330 768.345 929.850 771.175 ;
        RECT 5.330 762.905 929.850 765.735 ;
        RECT 5.330 757.465 929.850 760.295 ;
        RECT 5.330 752.025 929.850 754.855 ;
        RECT 5.330 746.585 929.850 749.415 ;
        RECT 5.330 741.145 929.850 743.975 ;
        RECT 5.330 735.705 929.850 738.535 ;
        RECT 5.330 730.265 929.850 733.095 ;
        RECT 5.330 724.825 929.850 727.655 ;
        RECT 5.330 719.385 929.850 722.215 ;
        RECT 5.330 713.945 929.850 716.775 ;
        RECT 5.330 708.505 929.850 711.335 ;
        RECT 5.330 703.065 929.850 705.895 ;
        RECT 5.330 697.625 929.850 700.455 ;
        RECT 5.330 692.185 929.850 695.015 ;
        RECT 5.330 686.745 929.850 689.575 ;
        RECT 5.330 681.305 929.850 684.135 ;
        RECT 5.330 675.865 929.850 678.695 ;
        RECT 5.330 670.425 929.850 673.255 ;
        RECT 5.330 664.985 929.850 667.815 ;
        RECT 5.330 659.545 929.850 662.375 ;
        RECT 5.330 654.105 929.850 656.935 ;
        RECT 5.330 648.665 929.850 651.495 ;
        RECT 5.330 643.225 929.850 646.055 ;
        RECT 5.330 637.785 929.850 640.615 ;
        RECT 5.330 632.345 929.850 635.175 ;
        RECT 5.330 626.905 929.850 629.735 ;
        RECT 5.330 621.465 929.850 624.295 ;
        RECT 5.330 616.025 929.850 618.855 ;
        RECT 5.330 610.585 929.850 613.415 ;
        RECT 5.330 605.145 929.850 607.975 ;
        RECT 5.330 599.705 929.850 602.535 ;
        RECT 5.330 594.265 929.850 597.095 ;
        RECT 5.330 588.825 929.850 591.655 ;
        RECT 5.330 583.385 929.850 586.215 ;
        RECT 5.330 577.945 929.850 580.775 ;
        RECT 5.330 572.505 929.850 575.335 ;
        RECT 5.330 567.065 929.850 569.895 ;
        RECT 5.330 561.625 929.850 564.455 ;
        RECT 5.330 556.185 929.850 559.015 ;
        RECT 5.330 550.745 929.850 553.575 ;
        RECT 5.330 545.305 929.850 548.135 ;
        RECT 5.330 539.865 929.850 542.695 ;
        RECT 5.330 534.425 929.850 537.255 ;
        RECT 5.330 528.985 929.850 531.815 ;
        RECT 5.330 523.545 929.850 526.375 ;
        RECT 5.330 518.105 929.850 520.935 ;
        RECT 5.330 512.665 929.850 515.495 ;
        RECT 5.330 507.225 929.850 510.055 ;
        RECT 5.330 501.785 929.850 504.615 ;
        RECT 5.330 496.345 929.850 499.175 ;
        RECT 5.330 490.905 929.850 493.735 ;
        RECT 5.330 485.465 929.850 488.295 ;
        RECT 5.330 480.025 929.850 482.855 ;
        RECT 5.330 474.585 929.850 477.415 ;
        RECT 5.330 469.145 929.850 471.975 ;
        RECT 5.330 463.705 929.850 466.535 ;
        RECT 5.330 458.265 929.850 461.095 ;
        RECT 5.330 452.825 929.850 455.655 ;
        RECT 5.330 447.385 929.850 450.215 ;
        RECT 5.330 441.945 929.850 444.775 ;
        RECT 5.330 436.505 929.850 439.335 ;
        RECT 5.330 431.065 929.850 433.895 ;
        RECT 5.330 425.625 929.850 428.455 ;
        RECT 5.330 420.185 929.850 423.015 ;
        RECT 5.330 414.745 929.850 417.575 ;
        RECT 5.330 409.305 929.850 412.135 ;
        RECT 5.330 403.865 929.850 406.695 ;
        RECT 5.330 398.425 929.850 401.255 ;
        RECT 5.330 392.985 929.850 395.815 ;
        RECT 5.330 387.545 929.850 390.375 ;
        RECT 5.330 382.105 929.850 384.935 ;
        RECT 5.330 376.665 929.850 379.495 ;
        RECT 5.330 371.225 929.850 374.055 ;
        RECT 5.330 365.785 929.850 368.615 ;
        RECT 5.330 360.345 929.850 363.175 ;
        RECT 5.330 354.905 929.850 357.735 ;
        RECT 5.330 349.465 929.850 352.295 ;
        RECT 5.330 344.025 929.850 346.855 ;
        RECT 5.330 338.585 929.850 341.415 ;
        RECT 5.330 333.145 929.850 335.975 ;
        RECT 5.330 327.705 929.850 330.535 ;
        RECT 5.330 322.265 929.850 325.095 ;
        RECT 5.330 316.825 929.850 319.655 ;
        RECT 5.330 311.385 929.850 314.215 ;
        RECT 5.330 305.945 929.850 308.775 ;
        RECT 5.330 300.505 929.850 303.335 ;
        RECT 5.330 295.065 929.850 297.895 ;
        RECT 5.330 289.625 929.850 292.455 ;
        RECT 5.330 284.185 929.850 287.015 ;
        RECT 5.330 278.745 929.850 281.575 ;
        RECT 5.330 273.305 929.850 276.135 ;
        RECT 5.330 267.865 929.850 270.695 ;
        RECT 5.330 262.425 929.850 265.255 ;
        RECT 5.330 256.985 929.850 259.815 ;
        RECT 5.330 251.545 929.850 254.375 ;
        RECT 5.330 246.105 929.850 248.935 ;
        RECT 5.330 240.665 929.850 243.495 ;
        RECT 5.330 235.225 929.850 238.055 ;
        RECT 5.330 229.785 929.850 232.615 ;
        RECT 5.330 224.345 929.850 227.175 ;
        RECT 5.330 218.905 929.850 221.735 ;
        RECT 5.330 213.465 929.850 216.295 ;
        RECT 5.330 208.025 929.850 210.855 ;
        RECT 5.330 202.585 929.850 205.415 ;
        RECT 5.330 197.145 929.850 199.975 ;
        RECT 5.330 191.705 929.850 194.535 ;
        RECT 5.330 186.265 929.850 189.095 ;
        RECT 5.330 180.825 929.850 183.655 ;
        RECT 5.330 175.385 929.850 178.215 ;
        RECT 5.330 169.945 929.850 172.775 ;
        RECT 5.330 164.505 929.850 167.335 ;
        RECT 5.330 159.065 929.850 161.895 ;
        RECT 5.330 153.625 929.850 156.455 ;
        RECT 5.330 148.185 929.850 151.015 ;
        RECT 5.330 142.745 929.850 145.575 ;
        RECT 5.330 137.305 929.850 140.135 ;
        RECT 5.330 131.865 929.850 134.695 ;
        RECT 5.330 126.425 929.850 129.255 ;
        RECT 5.330 120.985 929.850 123.815 ;
        RECT 5.330 115.545 929.850 118.375 ;
        RECT 5.330 110.105 929.850 112.935 ;
        RECT 5.330 104.665 929.850 107.495 ;
        RECT 5.330 99.225 929.850 102.055 ;
        RECT 5.330 93.785 929.850 96.615 ;
        RECT 5.330 88.345 929.850 91.175 ;
        RECT 5.330 82.905 929.850 85.735 ;
        RECT 5.330 77.465 929.850 80.295 ;
        RECT 5.330 72.025 929.850 74.855 ;
        RECT 5.330 66.585 929.850 69.415 ;
        RECT 5.330 61.145 929.850 63.975 ;
        RECT 5.330 55.705 929.850 58.535 ;
        RECT 5.330 50.265 929.850 53.095 ;
        RECT 5.330 44.825 929.850 47.655 ;
        RECT 5.330 39.385 929.850 42.215 ;
        RECT 5.330 33.945 929.850 36.775 ;
        RECT 5.330 28.505 929.850 31.335 ;
        RECT 5.330 23.065 929.850 25.895 ;
        RECT 5.330 17.625 929.850 20.455 ;
        RECT 5.330 12.185 929.850 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 929.660 933.045 ;
      LAYER met1 ;
        RECT 5.520 6.840 929.660 933.200 ;
      LAYER met2 ;
        RECT 7.450 4.280 927.660 933.145 ;
        RECT 8.010 3.670 18.670 4.280 ;
        RECT 19.510 3.670 30.170 4.280 ;
        RECT 31.010 3.670 41.670 4.280 ;
        RECT 42.510 3.670 53.170 4.280 ;
        RECT 54.010 3.670 64.670 4.280 ;
        RECT 65.510 3.670 76.170 4.280 ;
        RECT 77.010 3.670 87.670 4.280 ;
        RECT 88.510 3.670 99.170 4.280 ;
        RECT 100.010 3.670 110.670 4.280 ;
        RECT 111.510 3.670 122.170 4.280 ;
        RECT 123.010 3.670 133.670 4.280 ;
        RECT 134.510 3.670 145.170 4.280 ;
        RECT 146.010 3.670 156.670 4.280 ;
        RECT 157.510 3.670 168.170 4.280 ;
        RECT 169.010 3.670 179.670 4.280 ;
        RECT 180.510 3.670 191.170 4.280 ;
        RECT 192.010 3.670 202.670 4.280 ;
        RECT 203.510 3.670 214.170 4.280 ;
        RECT 215.010 3.670 225.670 4.280 ;
        RECT 226.510 3.670 237.170 4.280 ;
        RECT 238.010 3.670 248.670 4.280 ;
        RECT 249.510 3.670 260.170 4.280 ;
        RECT 261.010 3.670 271.670 4.280 ;
        RECT 272.510 3.670 283.170 4.280 ;
        RECT 284.010 3.670 294.670 4.280 ;
        RECT 295.510 3.670 306.170 4.280 ;
        RECT 307.010 3.670 317.670 4.280 ;
        RECT 318.510 3.670 329.170 4.280 ;
        RECT 330.010 3.670 340.670 4.280 ;
        RECT 341.510 3.670 352.170 4.280 ;
        RECT 353.010 3.670 363.670 4.280 ;
        RECT 364.510 3.670 375.170 4.280 ;
        RECT 376.010 3.670 386.670 4.280 ;
        RECT 387.510 3.670 398.170 4.280 ;
        RECT 399.010 3.670 409.670 4.280 ;
        RECT 410.510 3.670 421.170 4.280 ;
        RECT 422.010 3.670 432.670 4.280 ;
        RECT 433.510 3.670 444.170 4.280 ;
        RECT 445.010 3.670 455.670 4.280 ;
        RECT 456.510 3.670 467.170 4.280 ;
        RECT 468.010 3.670 478.670 4.280 ;
        RECT 479.510 3.670 490.170 4.280 ;
        RECT 491.010 3.670 501.670 4.280 ;
        RECT 502.510 3.670 513.170 4.280 ;
        RECT 514.010 3.670 524.670 4.280 ;
        RECT 525.510 3.670 536.170 4.280 ;
        RECT 537.010 3.670 547.670 4.280 ;
        RECT 548.510 3.670 559.170 4.280 ;
        RECT 560.010 3.670 570.670 4.280 ;
        RECT 571.510 3.670 582.170 4.280 ;
        RECT 583.010 3.670 593.670 4.280 ;
        RECT 594.510 3.670 605.170 4.280 ;
        RECT 606.010 3.670 616.670 4.280 ;
        RECT 617.510 3.670 628.170 4.280 ;
        RECT 629.010 3.670 639.670 4.280 ;
        RECT 640.510 3.670 651.170 4.280 ;
        RECT 652.010 3.670 662.670 4.280 ;
        RECT 663.510 3.670 674.170 4.280 ;
        RECT 675.010 3.670 685.670 4.280 ;
        RECT 686.510 3.670 697.170 4.280 ;
        RECT 698.010 3.670 708.670 4.280 ;
        RECT 709.510 3.670 720.170 4.280 ;
        RECT 721.010 3.670 731.670 4.280 ;
        RECT 732.510 3.670 743.170 4.280 ;
        RECT 744.010 3.670 754.670 4.280 ;
        RECT 755.510 3.670 766.170 4.280 ;
        RECT 767.010 3.670 777.670 4.280 ;
        RECT 778.510 3.670 789.170 4.280 ;
        RECT 790.010 3.670 800.670 4.280 ;
        RECT 801.510 3.670 812.170 4.280 ;
        RECT 813.010 3.670 823.670 4.280 ;
        RECT 824.510 3.670 835.170 4.280 ;
        RECT 836.010 3.670 846.670 4.280 ;
        RECT 847.510 3.670 858.170 4.280 ;
        RECT 859.010 3.670 869.670 4.280 ;
        RECT 870.510 3.670 881.170 4.280 ;
        RECT 882.010 3.670 892.670 4.280 ;
        RECT 893.510 3.670 904.170 4.280 ;
        RECT 905.010 3.670 915.670 4.280 ;
        RECT 916.510 3.670 927.170 4.280 ;
      LAYER met3 ;
        RECT 7.425 9.710 900.615 933.125 ;
      LAYER met4 ;
        RECT 15.015 10.375 20.640 858.665 ;
        RECT 23.040 10.375 97.440 858.665 ;
        RECT 99.840 10.375 174.240 858.665 ;
        RECT 176.640 10.375 251.040 858.665 ;
        RECT 253.440 10.375 327.840 858.665 ;
        RECT 330.240 10.375 404.640 858.665 ;
        RECT 407.040 10.375 481.440 858.665 ;
        RECT 483.840 10.375 558.240 858.665 ;
        RECT 560.640 10.375 635.040 858.665 ;
        RECT 637.440 10.375 711.840 858.665 ;
        RECT 714.240 10.375 788.640 858.665 ;
        RECT 791.040 10.375 865.440 858.665 ;
        RECT 867.840 10.375 895.785 858.665 ;
  END
END bec
END LIBRARY

