magic
tech sky130A
timestamp 1730450826
<< nwell >>
rect -130 -40 340 340
<< pwell >>
rect -130 -80 100 -70
rect 120 -80 340 -70
rect -130 -350 340 -80
<< nmos >>
rect 0 -310 120 -110
rect 160 -310 280 -110
<< pmos >>
rect 0 0 120 300
rect 160 0 280 300
<< ndiff >>
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -310 0 -300
rect 120 -120 160 -110
rect 120 -140 130 -120
rect 150 -140 160 -120
rect 120 -160 160 -140
rect 120 -180 130 -160
rect 150 -180 160 -160
rect 120 -200 160 -180
rect 120 -220 130 -200
rect 150 -220 160 -200
rect 120 -240 160 -220
rect 120 -260 130 -240
rect 150 -260 160 -240
rect 120 -280 160 -260
rect 120 -300 130 -280
rect 150 -300 160 -280
rect 120 -310 160 -300
rect 280 -120 320 -110
rect 280 -140 290 -120
rect 310 -140 320 -120
rect 280 -160 320 -140
rect 280 -180 290 -160
rect 310 -180 320 -160
rect 280 -200 320 -180
rect 280 -220 290 -200
rect 310 -220 320 -200
rect 280 -240 320 -220
rect 280 -260 290 -240
rect 310 -260 320 -240
rect 280 -280 320 -260
rect 280 -300 290 -280
rect 310 -300 320 -280
rect 280 -310 320 -300
<< pdiff >>
rect -40 290 0 300
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 120 290 160 300
rect 120 270 130 290
rect 150 270 160 290
rect 120 250 160 270
rect 120 230 130 250
rect 150 230 160 250
rect 120 210 160 230
rect 120 190 130 210
rect 150 190 160 210
rect 120 170 160 190
rect 120 150 130 170
rect 150 150 160 170
rect 120 130 160 150
rect 120 110 130 130
rect 150 110 160 130
rect 120 90 160 110
rect 120 70 130 90
rect 150 70 160 90
rect 120 50 160 70
rect 120 30 130 50
rect 150 30 160 50
rect 120 0 160 30
rect 280 290 320 300
rect 280 270 290 290
rect 310 270 320 290
rect 280 250 320 270
rect 280 230 290 250
rect 310 230 320 250
rect 280 210 320 230
rect 280 190 290 210
rect 310 190 320 210
rect 280 170 320 190
rect 280 150 290 170
rect 310 150 320 170
rect 280 130 320 150
rect 280 110 290 130
rect 310 110 320 130
rect 280 90 320 110
rect 280 70 290 90
rect 310 70 320 90
rect 280 50 320 70
rect 280 30 290 50
rect 310 30 320 50
rect 280 0 320 30
<< ndiffc >>
rect -30 -140 -10 -120
rect -30 -180 -10 -160
rect -30 -220 -10 -200
rect -30 -260 -10 -240
rect -30 -300 -10 -280
rect 130 -140 150 -120
rect 130 -180 150 -160
rect 130 -220 150 -200
rect 130 -260 150 -240
rect 130 -300 150 -280
rect 290 -140 310 -120
rect 290 -180 310 -160
rect 290 -220 310 -200
rect 290 -260 310 -240
rect 290 -300 310 -280
<< pdiffc >>
rect -30 270 -10 290
rect -30 230 -10 250
rect -30 190 -10 210
rect -30 150 -10 170
rect -30 110 -10 130
rect -30 70 -10 90
rect -30 30 -10 50
rect 130 270 150 290
rect 130 230 150 250
rect 130 190 150 210
rect 130 150 150 170
rect 130 110 150 130
rect 130 70 150 90
rect 130 30 150 50
rect 290 270 310 290
rect 290 230 310 250
rect 290 190 310 210
rect 290 150 310 170
rect 290 110 310 130
rect 290 70 310 90
rect 290 30 310 50
<< psubdiff >>
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< nsubdiff >>
rect -110 290 -70 305
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
<< psubdiffcont >>
rect -100 -300 -80 -280
<< nsubdiffcont >>
rect -100 270 -80 290
<< poly >>
rect 0 300 120 340
rect 160 300 280 340
rect 0 -40 120 0
rect 160 -40 280 0
rect 0 -45 280 -40
rect 0 -65 35 -45
rect 55 -65 200 -45
rect 220 -65 280 -45
rect 0 -70 280 -65
rect 0 -110 120 -70
rect 160 -110 280 -70
rect 0 -350 120 -310
rect 160 -350 280 -310
<< polycont >>
rect 35 -65 55 -45
rect 200 -65 220 -45
<< locali >>
rect -110 390 320 430
rect -110 290 -70 390
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
rect -40 290 0 390
rect -40 270 -30 290
rect -10 270 0 290
rect -40 250 0 270
rect -40 230 -30 250
rect -10 230 0 250
rect -40 210 0 230
rect -40 190 -30 210
rect -10 190 0 210
rect -40 170 0 190
rect -40 150 -30 170
rect -10 150 0 170
rect -40 130 0 150
rect -40 110 -30 130
rect -10 110 0 130
rect -40 90 0 110
rect -40 70 -30 90
rect -10 70 0 90
rect -40 50 0 70
rect -40 30 -30 50
rect -10 30 0 50
rect -40 0 0 30
rect 120 290 160 300
rect 120 270 130 290
rect 150 270 160 290
rect 120 250 160 270
rect 120 230 130 250
rect 150 230 160 250
rect 120 210 160 230
rect 120 190 130 210
rect 150 190 160 210
rect 120 170 160 190
rect 120 150 130 170
rect 150 150 160 170
rect 120 130 160 150
rect 120 110 130 130
rect 150 110 160 130
rect 120 90 160 110
rect 120 70 130 90
rect 150 70 160 90
rect 120 50 160 70
rect 120 30 130 50
rect 150 30 160 50
rect 25 -45 70 -35
rect 25 -65 35 -45
rect 55 -65 70 -45
rect 25 -80 70 -65
rect -40 -120 0 -110
rect -40 -140 -30 -120
rect -10 -140 0 -120
rect -40 -160 0 -140
rect -40 -180 -30 -160
rect -10 -180 0 -160
rect -40 -200 0 -180
rect -40 -220 -30 -200
rect -10 -220 0 -200
rect -40 -240 0 -220
rect -40 -260 -30 -240
rect -10 -260 0 -240
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -400 -70 -300
rect -40 -280 0 -260
rect -40 -300 -30 -280
rect -10 -300 0 -280
rect -40 -400 0 -300
rect 120 -120 160 30
rect 280 290 320 390
rect 280 270 290 290
rect 310 270 320 290
rect 280 250 320 270
rect 280 230 290 250
rect 310 230 320 250
rect 280 210 320 230
rect 280 190 290 210
rect 310 190 320 210
rect 280 170 320 190
rect 280 150 290 170
rect 310 150 320 170
rect 280 130 320 150
rect 280 110 290 130
rect 310 110 320 130
rect 280 90 320 110
rect 280 70 290 90
rect 310 70 320 90
rect 280 50 320 70
rect 280 30 290 50
rect 310 30 320 50
rect 280 0 320 30
rect 185 -45 230 -35
rect 185 -65 200 -45
rect 220 -65 230 -45
rect 185 -80 230 -65
rect 120 -140 130 -120
rect 150 -140 160 -120
rect 120 -160 160 -140
rect 120 -180 130 -160
rect 150 -180 160 -160
rect 120 -200 160 -180
rect 120 -220 130 -200
rect 150 -220 160 -200
rect 120 -240 160 -220
rect 120 -260 130 -240
rect 150 -260 160 -240
rect 120 -280 160 -260
rect 120 -300 130 -280
rect 150 -300 160 -280
rect 120 -310 160 -300
rect 280 -120 320 -110
rect 280 -140 290 -120
rect 310 -140 320 -120
rect 280 -160 320 -140
rect 280 -180 290 -160
rect 310 -180 320 -160
rect 280 -200 320 -180
rect 280 -220 290 -200
rect 310 -220 320 -200
rect 280 -240 320 -220
rect 280 -260 290 -240
rect 310 -260 320 -240
rect 280 -280 320 -260
rect 280 -300 290 -280
rect 310 -300 320 -280
rect 280 -400 320 -300
rect -110 -440 320 -400
<< viali >>
rect -100 270 -80 290
rect 35 -65 55 -45
rect -100 -300 -80 -280
rect 200 -65 220 -45
<< metal1 >>
rect -110 290 -70 305
rect -110 270 -100 290
rect -80 270 -70 290
rect -110 255 -70 270
rect 25 -45 230 -35
rect 25 -65 35 -45
rect 55 -65 200 -45
rect 220 -65 230 -45
rect 25 -80 230 -65
rect -110 -280 -70 -265
rect -110 -300 -100 -280
rect -80 -300 -70 -280
rect -110 -315 -70 -300
<< labels >>
rlabel metal1 25 -55 25 -55 7 A
port 1 w
rlabel locali -70 430 -70 430 1 VDDA
port 3 n
rlabel locali -70 -440 -70 -440 5 VGND
port 4 s
rlabel locali 140 -310 140 -310 5 Y
port 2 s
<< end >>
