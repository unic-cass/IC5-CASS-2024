magic
tech sky130A
magscale 1 2
timestamp 1731518408
<< nwell >>
rect 1066 104709 118902 105275
rect 1066 103621 118902 104187
rect 1066 102533 118902 103099
rect 1066 101445 118902 102011
rect 1066 100357 118902 100923
rect 1066 99269 118902 99835
rect 1066 98181 118902 98747
rect 1066 97093 118902 97659
rect 1066 96005 118902 96571
rect 1066 94917 118902 95483
rect 1066 93829 118902 94395
rect 1066 92741 118902 93307
rect 1066 91653 118902 92219
rect 1066 90565 118902 91131
rect 1066 89477 118902 90043
rect 1066 88389 118902 88955
rect 1066 87301 118902 87867
rect 1066 86213 118902 86779
rect 1066 85125 118902 85691
rect 1066 84037 118902 84603
rect 1066 82949 118902 83515
rect 1066 81861 118902 82427
rect 1066 80773 118902 81339
rect 1066 79685 118902 80251
rect 1066 78597 118902 79163
rect 1066 77509 118902 78075
rect 1066 76421 118902 76987
rect 1066 75333 118902 75899
rect 1066 74245 118902 74811
rect 1066 73157 118902 73723
rect 1066 72069 118902 72635
rect 1066 70981 118902 71547
rect 1066 69893 118902 70459
rect 1066 68805 118902 69371
rect 1066 67717 118902 68283
rect 1066 66629 118902 67195
rect 1066 65541 118902 66107
rect 1066 64453 118902 65019
rect 1066 63365 118902 63931
rect 1066 62277 118902 62843
rect 1066 61189 118902 61755
rect 1066 60101 118902 60667
rect 1066 59013 118902 59579
rect 1066 57925 118902 58491
rect 1066 56837 118902 57403
rect 1066 55749 118902 56315
rect 1066 54661 118902 55227
rect 1066 53573 118902 54139
rect 1066 52485 118902 53051
rect 1066 51397 118902 51963
rect 1066 50309 118902 50875
rect 1066 49221 118902 49787
rect 1066 48133 118902 48699
rect 1066 47045 118902 47611
rect 1066 45957 118902 46523
rect 1066 44869 118902 45435
rect 1066 43781 118902 44347
rect 1066 42693 118902 43259
rect 1066 41605 118902 42171
rect 1066 40517 118902 41083
rect 1066 39429 118902 39995
rect 1066 38341 118902 38907
rect 1066 37253 118902 37819
rect 1066 36165 118902 36731
rect 1066 35077 118902 35643
rect 1066 33989 118902 34555
rect 1066 32901 118902 33467
rect 1066 31813 118902 32379
rect 1066 30725 118902 31291
rect 1066 29637 118902 30203
rect 1066 28549 118902 29115
rect 1066 27461 118902 28027
rect 1066 26373 118902 26939
rect 1066 25285 118902 25851
rect 1066 24197 118902 24763
rect 1066 23109 118902 23675
rect 1066 22021 118902 22587
rect 1066 20933 118902 21499
rect 1066 19845 118902 20411
rect 1066 18757 118902 19323
rect 1066 17669 118902 18235
rect 1066 16581 118902 17147
rect 1066 15493 118902 16059
rect 1066 14405 118902 14971
rect 1066 13317 118902 13883
rect 1066 12229 118902 12795
rect 1066 11141 118902 11707
rect 1066 10053 118902 10619
rect 1066 8965 118902 9531
rect 1066 7877 118902 8443
rect 1066 6789 118902 7355
rect 1066 5701 118902 6267
rect 1066 4613 118902 5179
rect 1066 3525 118902 4091
rect 1066 2437 118902 3003
<< obsli1 >>
rect 1104 2159 118864 105553
<< obsm1 >>
rect 1104 2128 118942 105584
<< metal2 >>
rect 6090 107200 6146 108000
rect 18050 107200 18106 108000
rect 30010 107200 30066 108000
rect 41970 107200 42026 108000
rect 53930 107200 53986 108000
rect 65890 107200 65946 108000
rect 77850 107200 77906 108000
rect 89810 107200 89866 108000
rect 101770 107200 101826 108000
rect 113730 107200 113786 108000
<< obsm2 >>
rect 3976 107144 6034 107200
rect 6202 107144 17994 107200
rect 18162 107144 29954 107200
rect 30122 107144 41914 107200
rect 42082 107144 53874 107200
rect 54042 107144 65834 107200
rect 66002 107144 77794 107200
rect 77962 107144 89754 107200
rect 89922 107144 101714 107200
rect 101882 107144 113674 107200
rect 113842 107144 118938 107200
rect 3976 2139 118938 107144
<< metal3 >>
rect 119200 103096 120000 103216
rect 119200 94120 120000 94240
rect 119200 85144 120000 85264
rect 119200 76168 120000 76288
rect 119200 67192 120000 67312
rect 119200 58216 120000 58336
rect 119200 49240 120000 49360
rect 119200 40264 120000 40384
rect 119200 31288 120000 31408
rect 119200 22312 120000 22432
rect 119200 13336 120000 13456
rect 119200 4360 120000 4480
<< obsm3 >>
rect 4210 103296 119200 105569
rect 4210 103016 119120 103296
rect 4210 94320 119200 103016
rect 4210 94040 119120 94320
rect 4210 85344 119200 94040
rect 4210 85064 119120 85344
rect 4210 76368 119200 85064
rect 4210 76088 119120 76368
rect 4210 67392 119200 76088
rect 4210 67112 119120 67392
rect 4210 58416 119200 67112
rect 4210 58136 119120 58416
rect 4210 49440 119200 58136
rect 4210 49160 119120 49440
rect 4210 40464 119200 49160
rect 4210 40184 119120 40464
rect 4210 31488 119200 40184
rect 4210 31208 119120 31488
rect 4210 22512 119200 31208
rect 4210 22232 119120 22512
rect 4210 13536 119200 22232
rect 4210 13256 119120 13536
rect 4210 4560 119200 13256
rect 4210 4280 119120 4560
rect 4210 2143 119200 4280
<< metal4 >>
rect 4208 2128 4528 105584
rect 19568 2128 19888 105584
rect 34928 2128 35248 105584
rect 50288 2128 50608 105584
rect 65648 2128 65968 105584
rect 81008 2128 81328 105584
rect 96368 2128 96688 105584
rect 111728 2128 112048 105584
<< obsm4 >>
rect 14411 7379 19488 99925
rect 19968 7379 34848 99925
rect 35328 7379 50208 99925
rect 50688 7379 65568 99925
rect 66048 7379 80928 99925
rect 81408 7379 96288 99925
rect 96768 7379 111648 99925
rect 112128 7379 115677 99925
<< obsm5 >>
rect 24588 34180 84340 68500
<< labels >>
rlabel metal2 s 89810 107200 89866 108000 6 clk
port 1 nsew signal input
rlabel metal3 s 119200 103096 120000 103216 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 119200 85144 120000 85264 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 119200 67192 120000 67312 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 119200 49240 120000 49360 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 119200 31288 120000 31408 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 119200 13336 120000 13456 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 53930 107200 53986 108000 6 io_oeb[0]
port 8 nsew signal output
rlabel metal2 s 77850 107200 77906 108000 6 io_oeb[10]
port 9 nsew signal output
rlabel metal2 s 30010 107200 30066 108000 6 io_oeb[1]
port 10 nsew signal output
rlabel metal2 s 6090 107200 6146 108000 6 io_oeb[2]
port 11 nsew signal output
rlabel metal3 s 119200 94120 120000 94240 6 io_oeb[3]
port 12 nsew signal output
rlabel metal3 s 119200 76168 120000 76288 6 io_oeb[4]
port 13 nsew signal output
rlabel metal3 s 119200 58216 120000 58336 6 io_oeb[5]
port 14 nsew signal output
rlabel metal3 s 119200 40264 120000 40384 6 io_oeb[6]
port 15 nsew signal output
rlabel metal3 s 119200 22312 120000 22432 6 io_oeb[7]
port 16 nsew signal output
rlabel metal3 s 119200 4360 120000 4480 6 io_oeb[8]
port 17 nsew signal output
rlabel metal2 s 101770 107200 101826 108000 6 io_oeb[9]
port 18 nsew signal output
rlabel metal2 s 65890 107200 65946 108000 6 io_out[0]
port 19 nsew signal output
rlabel metal2 s 41970 107200 42026 108000 6 io_out[1]
port 20 nsew signal output
rlabel metal2 s 18050 107200 18106 108000 6 io_out[2]
port 21 nsew signal output
rlabel metal2 s 113730 107200 113786 108000 6 rst
port 22 nsew signal input
rlabel metal4 s 4208 2128 4528 105584 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 105584 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 105584 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 105584 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 105584 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 105584 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 105584 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 105584 6 vssd1
port 24 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 108000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36111658
string GDS_FILE /home/cass/projects/IC5-CASS-2024/openlane/hs_ascon/runs/24_11_13_23_52/results/signoff/ascon_wrapper.magic.gds
string GDS_START 844014
<< end >>

