magic
tech sky130A
magscale 1 2
timestamp 1731168528
<< nwell >>
rect 1066 251589 251750 252155
rect 1066 250501 251750 251067
rect 1066 249413 251750 249979
rect 1066 248325 251750 248891
rect 1066 247237 251750 247803
rect 1066 246149 251750 246715
rect 1066 245061 251750 245627
rect 1066 243973 251750 244539
rect 1066 242885 251750 243451
rect 1066 241797 251750 242363
rect 1066 240709 251750 241275
rect 1066 239621 251750 240187
rect 1066 238533 251750 239099
rect 1066 237445 251750 238011
rect 1066 236357 251750 236923
rect 1066 235269 251750 235835
rect 1066 234181 251750 234747
rect 1066 233093 251750 233659
rect 1066 232005 251750 232571
rect 1066 230917 251750 231483
rect 1066 229829 251750 230395
rect 1066 228741 251750 229307
rect 1066 227653 251750 228219
rect 1066 226565 251750 227131
rect 1066 225477 251750 226043
rect 1066 224389 251750 224955
rect 1066 223301 251750 223867
rect 1066 222213 251750 222779
rect 1066 221125 251750 221691
rect 1066 220037 251750 220603
rect 1066 218949 251750 219515
rect 1066 217861 251750 218427
rect 1066 216773 251750 217339
rect 1066 215685 251750 216251
rect 1066 214597 251750 215163
rect 1066 213509 251750 214075
rect 1066 212421 251750 212987
rect 1066 211333 251750 211899
rect 1066 210245 251750 210811
rect 1066 209157 251750 209723
rect 1066 208069 251750 208635
rect 1066 206981 251750 207547
rect 1066 205893 251750 206459
rect 1066 204805 251750 205371
rect 1066 203717 251750 204283
rect 1066 202629 251750 203195
rect 1066 201541 251750 202107
rect 1066 200453 251750 201019
rect 1066 199365 251750 199931
rect 1066 198277 251750 198843
rect 1066 197189 251750 197755
rect 1066 196101 251750 196667
rect 1066 195013 251750 195579
rect 1066 193925 251750 194491
rect 1066 192837 251750 193403
rect 1066 191749 251750 192315
rect 1066 190661 251750 191227
rect 1066 189573 251750 190139
rect 1066 188485 251750 189051
rect 1066 187397 251750 187963
rect 1066 186309 251750 186875
rect 1066 185221 251750 185787
rect 1066 184133 251750 184699
rect 1066 183045 251750 183611
rect 1066 181957 251750 182523
rect 1066 180869 251750 181435
rect 1066 179781 251750 180347
rect 1066 178693 251750 179259
rect 1066 177605 251750 178171
rect 1066 176517 251750 177083
rect 1066 175429 251750 175995
rect 1066 174341 251750 174907
rect 1066 173253 251750 173819
rect 1066 172165 251750 172731
rect 1066 171077 251750 171643
rect 1066 169989 251750 170555
rect 1066 168901 251750 169467
rect 1066 167813 251750 168379
rect 1066 166725 251750 167291
rect 1066 165637 251750 166203
rect 1066 164549 251750 165115
rect 1066 163461 251750 164027
rect 1066 162373 251750 162939
rect 1066 161285 251750 161851
rect 1066 160197 251750 160763
rect 1066 159109 251750 159675
rect 1066 158021 251750 158587
rect 1066 156933 251750 157499
rect 1066 155845 251750 156411
rect 1066 154757 251750 155323
rect 1066 153669 251750 154235
rect 1066 152581 251750 153147
rect 1066 151493 251750 152059
rect 1066 150405 251750 150971
rect 1066 149317 251750 149883
rect 1066 148229 251750 148795
rect 1066 147141 251750 147707
rect 1066 146053 251750 146619
rect 1066 144965 251750 145531
rect 1066 143877 251750 144443
rect 1066 142789 251750 143355
rect 1066 141701 251750 142267
rect 1066 140613 251750 141179
rect 1066 139525 251750 140091
rect 1066 138437 251750 139003
rect 1066 137349 251750 137915
rect 1066 136261 251750 136827
rect 1066 135173 251750 135739
rect 1066 134085 251750 134651
rect 1066 132997 251750 133563
rect 1066 131909 251750 132475
rect 1066 130821 251750 131387
rect 1066 129733 251750 130299
rect 1066 128645 251750 129211
rect 1066 127557 251750 128123
rect 1066 126469 251750 127035
rect 1066 125381 251750 125947
rect 1066 124293 251750 124859
rect 1066 123205 251750 123771
rect 1066 122117 251750 122683
rect 1066 121029 251750 121595
rect 1066 119941 251750 120507
rect 1066 118853 251750 119419
rect 1066 117765 251750 118331
rect 1066 116677 251750 117243
rect 1066 115589 251750 116155
rect 1066 114501 251750 115067
rect 1066 113413 251750 113979
rect 1066 112325 251750 112891
rect 1066 111237 251750 111803
rect 1066 110149 251750 110715
rect 1066 109061 251750 109627
rect 1066 107973 251750 108539
rect 1066 106885 251750 107451
rect 1066 105797 251750 106363
rect 1066 104709 251750 105275
rect 1066 103621 251750 104187
rect 1066 102533 251750 103099
rect 1066 101445 251750 102011
rect 1066 100357 251750 100923
rect 1066 99269 251750 99835
rect 1066 98181 251750 98747
rect 1066 97093 251750 97659
rect 1066 96005 251750 96571
rect 1066 94917 251750 95483
rect 1066 93829 251750 94395
rect 1066 92741 251750 93307
rect 1066 91653 251750 92219
rect 1066 90565 251750 91131
rect 1066 89477 251750 90043
rect 1066 88389 251750 88955
rect 1066 87301 251750 87867
rect 1066 86213 251750 86779
rect 1066 85125 251750 85691
rect 1066 84037 251750 84603
rect 1066 82949 251750 83515
rect 1066 81861 251750 82427
rect 1066 80773 251750 81339
rect 1066 79685 251750 80251
rect 1066 78597 251750 79163
rect 1066 77509 251750 78075
rect 1066 76421 251750 76987
rect 1066 75333 251750 75899
rect 1066 74245 251750 74811
rect 1066 73157 251750 73723
rect 1066 72069 251750 72635
rect 1066 70981 251750 71547
rect 1066 69893 251750 70459
rect 1066 68805 251750 69371
rect 1066 67717 251750 68283
rect 1066 66629 251750 67195
rect 1066 65541 251750 66107
rect 1066 64453 251750 65019
rect 1066 63365 251750 63931
rect 1066 62277 251750 62843
rect 1066 61189 251750 61755
rect 1066 60101 251750 60667
rect 1066 59013 251750 59579
rect 1066 57925 251750 58491
rect 1066 56837 251750 57403
rect 1066 55749 251750 56315
rect 1066 54661 251750 55227
rect 1066 53573 251750 54139
rect 1066 52485 251750 53051
rect 1066 51397 251750 51963
rect 1066 50309 251750 50875
rect 1066 49221 251750 49787
rect 1066 48133 251750 48699
rect 1066 47045 251750 47611
rect 1066 45957 251750 46523
rect 1066 44869 251750 45435
rect 1066 43781 251750 44347
rect 1066 42693 251750 43259
rect 1066 41605 251750 42171
rect 1066 40517 251750 41083
rect 1066 39429 251750 39995
rect 1066 38341 251750 38907
rect 1066 37253 251750 37819
rect 1066 36165 251750 36731
rect 1066 35077 251750 35643
rect 1066 33989 251750 34555
rect 1066 32901 251750 33467
rect 1066 31813 251750 32379
rect 1066 30725 251750 31291
rect 1066 29637 251750 30203
rect 1066 28549 251750 29115
rect 1066 27461 251750 28027
rect 1066 26373 251750 26939
rect 1066 25285 251750 25851
rect 1066 24197 251750 24763
rect 1066 23109 251750 23675
rect 1066 22021 251750 22587
rect 1066 20933 251750 21499
rect 1066 19845 251750 20411
rect 1066 18757 251750 19323
rect 1066 17669 251750 18235
rect 1066 16581 251750 17147
rect 1066 15493 251750 16059
rect 1066 14405 251750 14971
rect 1066 13317 251750 13883
rect 1066 12229 251750 12795
rect 1066 11141 251750 11707
rect 1066 10053 251750 10619
rect 1066 8965 251750 9531
rect 1066 7877 251750 8443
rect 1066 6789 251750 7355
rect 1066 5701 251750 6267
rect 1066 4613 251750 5179
rect 1066 3525 251750 4091
rect 1066 2437 251750 3003
<< obsli1 >>
rect 1104 2159 251712 252433
<< obsm1 >>
rect 1104 1096 252434 252464
<< metal2 >>
rect 63222 254232 63278 255032
rect 189630 254232 189686 255032
rect 5630 0 5686 800
rect 7930 0 7986 800
rect 10230 0 10286 800
rect 12530 0 12586 800
rect 14830 0 14886 800
rect 17130 0 17186 800
rect 19430 0 19486 800
rect 21730 0 21786 800
rect 24030 0 24086 800
rect 26330 0 26386 800
rect 28630 0 28686 800
rect 30930 0 30986 800
rect 33230 0 33286 800
rect 35530 0 35586 800
rect 37830 0 37886 800
rect 40130 0 40186 800
rect 42430 0 42486 800
rect 44730 0 44786 800
rect 47030 0 47086 800
rect 49330 0 49386 800
rect 51630 0 51686 800
rect 53930 0 53986 800
rect 56230 0 56286 800
rect 58530 0 58586 800
rect 60830 0 60886 800
rect 63130 0 63186 800
rect 65430 0 65486 800
rect 67730 0 67786 800
rect 70030 0 70086 800
rect 72330 0 72386 800
rect 74630 0 74686 800
rect 76930 0 76986 800
rect 79230 0 79286 800
rect 81530 0 81586 800
rect 83830 0 83886 800
rect 86130 0 86186 800
rect 88430 0 88486 800
rect 90730 0 90786 800
rect 93030 0 93086 800
rect 95330 0 95386 800
rect 97630 0 97686 800
rect 99930 0 99986 800
rect 102230 0 102286 800
rect 104530 0 104586 800
rect 106830 0 106886 800
rect 109130 0 109186 800
rect 111430 0 111486 800
rect 113730 0 113786 800
rect 116030 0 116086 800
rect 118330 0 118386 800
rect 120630 0 120686 800
rect 122930 0 122986 800
rect 125230 0 125286 800
rect 127530 0 127586 800
rect 129830 0 129886 800
rect 132130 0 132186 800
rect 134430 0 134486 800
rect 136730 0 136786 800
rect 139030 0 139086 800
rect 141330 0 141386 800
rect 143630 0 143686 800
rect 145930 0 145986 800
rect 148230 0 148286 800
rect 150530 0 150586 800
rect 152830 0 152886 800
rect 155130 0 155186 800
rect 157430 0 157486 800
rect 159730 0 159786 800
rect 162030 0 162086 800
rect 164330 0 164386 800
rect 166630 0 166686 800
rect 168930 0 168986 800
rect 171230 0 171286 800
rect 173530 0 173586 800
rect 175830 0 175886 800
rect 178130 0 178186 800
rect 180430 0 180486 800
rect 182730 0 182786 800
rect 185030 0 185086 800
rect 187330 0 187386 800
rect 189630 0 189686 800
rect 191930 0 191986 800
rect 194230 0 194286 800
rect 196530 0 196586 800
rect 198830 0 198886 800
rect 201130 0 201186 800
rect 203430 0 203486 800
rect 205730 0 205786 800
rect 208030 0 208086 800
rect 210330 0 210386 800
rect 212630 0 212686 800
rect 214930 0 214986 800
rect 217230 0 217286 800
rect 219530 0 219586 800
rect 221830 0 221886 800
rect 224130 0 224186 800
rect 226430 0 226486 800
rect 228730 0 228786 800
rect 231030 0 231086 800
rect 233330 0 233386 800
rect 235630 0 235686 800
rect 237930 0 237986 800
rect 240230 0 240286 800
rect 242530 0 242586 800
rect 244830 0 244886 800
rect 247130 0 247186 800
<< obsm2 >>
rect 2228 254176 63166 254232
rect 63334 254176 189574 254232
rect 189742 254176 252428 254232
rect 2228 856 252428 254176
rect 2228 734 5574 856
rect 5742 734 7874 856
rect 8042 734 10174 856
rect 10342 734 12474 856
rect 12642 734 14774 856
rect 14942 734 17074 856
rect 17242 734 19374 856
rect 19542 734 21674 856
rect 21842 734 23974 856
rect 24142 734 26274 856
rect 26442 734 28574 856
rect 28742 734 30874 856
rect 31042 734 33174 856
rect 33342 734 35474 856
rect 35642 734 37774 856
rect 37942 734 40074 856
rect 40242 734 42374 856
rect 42542 734 44674 856
rect 44842 734 46974 856
rect 47142 734 49274 856
rect 49442 734 51574 856
rect 51742 734 53874 856
rect 54042 734 56174 856
rect 56342 734 58474 856
rect 58642 734 60774 856
rect 60942 734 63074 856
rect 63242 734 65374 856
rect 65542 734 67674 856
rect 67842 734 69974 856
rect 70142 734 72274 856
rect 72442 734 74574 856
rect 74742 734 76874 856
rect 77042 734 79174 856
rect 79342 734 81474 856
rect 81642 734 83774 856
rect 83942 734 86074 856
rect 86242 734 88374 856
rect 88542 734 90674 856
rect 90842 734 92974 856
rect 93142 734 95274 856
rect 95442 734 97574 856
rect 97742 734 99874 856
rect 100042 734 102174 856
rect 102342 734 104474 856
rect 104642 734 106774 856
rect 106942 734 109074 856
rect 109242 734 111374 856
rect 111542 734 113674 856
rect 113842 734 115974 856
rect 116142 734 118274 856
rect 118442 734 120574 856
rect 120742 734 122874 856
rect 123042 734 125174 856
rect 125342 734 127474 856
rect 127642 734 129774 856
rect 129942 734 132074 856
rect 132242 734 134374 856
rect 134542 734 136674 856
rect 136842 734 138974 856
rect 139142 734 141274 856
rect 141442 734 143574 856
rect 143742 734 145874 856
rect 146042 734 148174 856
rect 148342 734 150474 856
rect 150642 734 152774 856
rect 152942 734 155074 856
rect 155242 734 157374 856
rect 157542 734 159674 856
rect 159842 734 161974 856
rect 162142 734 164274 856
rect 164442 734 166574 856
rect 166742 734 168874 856
rect 169042 734 171174 856
rect 171342 734 173474 856
rect 173642 734 175774 856
rect 175942 734 178074 856
rect 178242 734 180374 856
rect 180542 734 182674 856
rect 182842 734 184974 856
rect 185142 734 187274 856
rect 187442 734 189574 856
rect 189742 734 191874 856
rect 192042 734 194174 856
rect 194342 734 196474 856
rect 196642 734 198774 856
rect 198942 734 201074 856
rect 201242 734 203374 856
rect 203542 734 205674 856
rect 205842 734 207974 856
rect 208142 734 210274 856
rect 210442 734 212574 856
rect 212742 734 214874 856
rect 215042 734 217174 856
rect 217342 734 219474 856
rect 219642 734 221774 856
rect 221942 734 224074 856
rect 224242 734 226374 856
rect 226542 734 228674 856
rect 228842 734 230974 856
rect 231142 734 233274 856
rect 233442 734 235574 856
rect 235742 734 237874 856
rect 238042 734 240174 856
rect 240342 734 242474 856
rect 242642 734 244774 856
rect 244942 734 247074 856
rect 247242 734 252428 856
<< obsm3 >>
rect 4210 1667 250779 252449
<< metal4 >>
rect 4208 2128 4528 252464
rect 19568 2128 19888 252464
rect 34928 2128 35248 252464
rect 50288 2128 50608 252464
rect 65648 2128 65968 252464
rect 81008 2128 81328 252464
rect 96368 2128 96688 252464
rect 111728 2128 112048 252464
rect 127088 2128 127408 252464
rect 142448 2128 142768 252464
rect 157808 2128 158128 252464
rect 173168 2128 173488 252464
rect 188528 2128 188848 252464
rect 203888 2128 204208 252464
rect 219248 2128 219568 252464
rect 234608 2128 234928 252464
rect 249968 2128 250288 252464
<< obsm4 >>
rect 5027 3979 19488 252245
rect 19968 3979 34848 252245
rect 35328 3979 50208 252245
rect 50688 3979 65568 252245
rect 66048 3979 80928 252245
rect 81408 3979 96288 252245
rect 96768 3979 111648 252245
rect 112128 3979 127008 252245
rect 127488 3979 142368 252245
rect 142848 3979 157728 252245
rect 158208 3979 173088 252245
rect 173568 3979 188448 252245
rect 188928 3979 203808 252245
rect 204288 3979 219168 252245
rect 219648 3979 234528 252245
rect 235008 3979 249888 252245
rect 250368 3979 250733 252245
<< labels >>
rlabel metal2 s 63222 254232 63278 255032 6 phase_in
port 1 nsew signal input
rlabel metal4 s 4208 2128 4528 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 252464 6 vccd1
port 2 nsew power bidirectional
rlabel metal2 s 189630 254232 189686 255032 6 vco_enb_o
port 3 nsew signal output
rlabel metal4 s 19568 2128 19888 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 252464 6 vssd1
port 4 nsew ground bidirectional
rlabel metal2 s 5630 0 5686 800 6 wb_clk_i
port 5 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wb_rst_i
port 6 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_ack_o
port 7 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[0]
port 8 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_adr_i[10]
port 9 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 wbs_adr_i[11]
port 10 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 wbs_adr_i[12]
port 11 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 wbs_adr_i[13]
port 12 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 wbs_adr_i[14]
port 13 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 wbs_adr_i[15]
port 14 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 wbs_adr_i[16]
port 15 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 wbs_adr_i[17]
port 16 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 wbs_adr_i[18]
port 17 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 wbs_adr_i[19]
port 18 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[1]
port 19 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 wbs_adr_i[20]
port 20 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 wbs_adr_i[21]
port 21 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 wbs_adr_i[22]
port 22 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 wbs_adr_i[23]
port 23 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 wbs_adr_i[24]
port 24 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 wbs_adr_i[25]
port 25 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 wbs_adr_i[26]
port 26 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 wbs_adr_i[27]
port 27 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 wbs_adr_i[28]
port 28 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 wbs_adr_i[29]
port 29 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[2]
port 30 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 wbs_adr_i[30]
port 31 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 wbs_adr_i[31]
port 32 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[3]
port 33 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[4]
port 34 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wbs_adr_i[5]
port 35 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_adr_i[6]
port 36 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[7]
port 37 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wbs_adr_i[8]
port 38 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 wbs_adr_i[9]
port 39 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_cyc_i
port 40 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[0]
port 41 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_i[10]
port 42 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 wbs_dat_i[11]
port 43 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wbs_dat_i[12]
port 44 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 wbs_dat_i[13]
port 45 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 wbs_dat_i[14]
port 46 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 wbs_dat_i[15]
port 47 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 wbs_dat_i[16]
port 48 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 wbs_dat_i[17]
port 49 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 wbs_dat_i[18]
port 50 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 wbs_dat_i[19]
port 51 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[1]
port 52 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 wbs_dat_i[20]
port 53 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 wbs_dat_i[21]
port 54 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 wbs_dat_i[22]
port 55 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 wbs_dat_i[23]
port 56 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 wbs_dat_i[24]
port 57 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 wbs_dat_i[25]
port 58 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 wbs_dat_i[26]
port 59 nsew signal input
rlabel metal2 s 217230 0 217286 800 6 wbs_dat_i[27]
port 60 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 wbs_dat_i[28]
port 61 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 wbs_dat_i[29]
port 62 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[2]
port 63 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 wbs_dat_i[30]
port 64 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 wbs_dat_i[31]
port 65 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_i[3]
port 66 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_i[4]
port 67 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_dat_i[5]
port 68 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 wbs_dat_i[6]
port 69 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_dat_i[7]
port 70 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 wbs_dat_i[8]
port 71 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 wbs_dat_i[9]
port 72 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[0]
port 73 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 wbs_dat_o[10]
port 74 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 wbs_dat_o[11]
port 75 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[12]
port 76 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 wbs_dat_o[13]
port 77 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 wbs_dat_o[14]
port 78 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 wbs_dat_o[15]
port 79 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 wbs_dat_o[16]
port 80 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 wbs_dat_o[17]
port 81 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 wbs_dat_o[18]
port 82 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 wbs_dat_o[19]
port 83 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[1]
port 84 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 wbs_dat_o[20]
port 85 nsew signal output
rlabel metal2 s 178130 0 178186 800 6 wbs_dat_o[21]
port 86 nsew signal output
rlabel metal2 s 185030 0 185086 800 6 wbs_dat_o[22]
port 87 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 wbs_dat_o[23]
port 88 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 wbs_dat_o[24]
port 89 nsew signal output
rlabel metal2 s 205730 0 205786 800 6 wbs_dat_o[25]
port 90 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 wbs_dat_o[26]
port 91 nsew signal output
rlabel metal2 s 219530 0 219586 800 6 wbs_dat_o[27]
port 92 nsew signal output
rlabel metal2 s 226430 0 226486 800 6 wbs_dat_o[28]
port 93 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 wbs_dat_o[29]
port 94 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_o[2]
port 95 nsew signal output
rlabel metal2 s 240230 0 240286 800 6 wbs_dat_o[30]
port 96 nsew signal output
rlabel metal2 s 247130 0 247186 800 6 wbs_dat_o[31]
port 97 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[3]
port 98 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_o[4]
port 99 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 wbs_dat_o[5]
port 100 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_o[6]
port 101 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[7]
port 102 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 wbs_dat_o[8]
port 103 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_o[9]
port 104 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_sel_i[0]
port 105 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_sel_i[1]
port 106 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_sel_i[2]
port 107 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_sel_i[3]
port 108 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_stb_i
port 109 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_we_i
port 110 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 252888 255032
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 193154144
string GDS_FILE /home/admin/projects/IC5-CASS-2024_2/openlane/vco_adc_wrapper/runs/24_11_09_20_32/results/signoff/vco_adc_wrapper.magic.gds
string GDS_START 1077234
<< end >>

