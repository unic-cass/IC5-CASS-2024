VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bec
  CLASS BLOCK ;
  FOREIGN bec ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 650.000 ;
  PIN becStatus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END becStatus[0]
  PIN becStatus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END becStatus[1]
  PIN becStatus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END becStatus[2]
  PIN becStatus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END becStatus[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END data_out[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END enable
  PIN ki
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END ki
  PIN load_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END load_data
  PIN load_status[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END load_status[0]
  PIN load_status[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END load_status[1]
  PIN load_status[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END load_status[2]
  PIN load_status[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END load_status[3]
  PIN load_status[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END load_status[4]
  PIN load_status[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END load_status[5]
  PIN next_key
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END next_key
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END rst
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 636.720 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 636.720 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 636.565 ;
      LAYER met1 ;
        RECT 0.990 0.380 799.410 636.720 ;
      LAYER met2 ;
        RECT 1.020 4.280 799.380 636.665 ;
        RECT 1.020 0.155 13.150 4.280 ;
        RECT 13.990 0.155 22.810 4.280 ;
        RECT 23.650 0.155 32.470 4.280 ;
        RECT 33.310 0.155 42.130 4.280 ;
        RECT 42.970 0.155 51.790 4.280 ;
        RECT 52.630 0.155 61.450 4.280 ;
        RECT 62.290 0.155 71.110 4.280 ;
        RECT 71.950 0.155 80.770 4.280 ;
        RECT 81.610 0.155 90.430 4.280 ;
        RECT 91.270 0.155 100.090 4.280 ;
        RECT 100.930 0.155 109.750 4.280 ;
        RECT 110.590 0.155 119.410 4.280 ;
        RECT 120.250 0.155 129.070 4.280 ;
        RECT 129.910 0.155 138.730 4.280 ;
        RECT 139.570 0.155 148.390 4.280 ;
        RECT 149.230 0.155 158.050 4.280 ;
        RECT 158.890 0.155 167.710 4.280 ;
        RECT 168.550 0.155 177.370 4.280 ;
        RECT 178.210 0.155 187.030 4.280 ;
        RECT 187.870 0.155 196.690 4.280 ;
        RECT 197.530 0.155 206.350 4.280 ;
        RECT 207.190 0.155 216.010 4.280 ;
        RECT 216.850 0.155 225.670 4.280 ;
        RECT 226.510 0.155 235.330 4.280 ;
        RECT 236.170 0.155 244.990 4.280 ;
        RECT 245.830 0.155 254.650 4.280 ;
        RECT 255.490 0.155 264.310 4.280 ;
        RECT 265.150 0.155 273.970 4.280 ;
        RECT 274.810 0.155 283.630 4.280 ;
        RECT 284.470 0.155 293.290 4.280 ;
        RECT 294.130 0.155 302.950 4.280 ;
        RECT 303.790 0.155 312.610 4.280 ;
        RECT 313.450 0.155 322.270 4.280 ;
        RECT 323.110 0.155 331.930 4.280 ;
        RECT 332.770 0.155 341.590 4.280 ;
        RECT 342.430 0.155 351.250 4.280 ;
        RECT 352.090 0.155 360.910 4.280 ;
        RECT 361.750 0.155 370.570 4.280 ;
        RECT 371.410 0.155 380.230 4.280 ;
        RECT 381.070 0.155 389.890 4.280 ;
        RECT 390.730 0.155 399.550 4.280 ;
        RECT 400.390 0.155 409.210 4.280 ;
        RECT 410.050 0.155 418.870 4.280 ;
        RECT 419.710 0.155 428.530 4.280 ;
        RECT 429.370 0.155 438.190 4.280 ;
        RECT 439.030 0.155 447.850 4.280 ;
        RECT 448.690 0.155 457.510 4.280 ;
        RECT 458.350 0.155 467.170 4.280 ;
        RECT 468.010 0.155 476.830 4.280 ;
        RECT 477.670 0.155 486.490 4.280 ;
        RECT 487.330 0.155 496.150 4.280 ;
        RECT 496.990 0.155 505.810 4.280 ;
        RECT 506.650 0.155 515.470 4.280 ;
        RECT 516.310 0.155 525.130 4.280 ;
        RECT 525.970 0.155 534.790 4.280 ;
        RECT 535.630 0.155 544.450 4.280 ;
        RECT 545.290 0.155 554.110 4.280 ;
        RECT 554.950 0.155 563.770 4.280 ;
        RECT 564.610 0.155 573.430 4.280 ;
        RECT 574.270 0.155 583.090 4.280 ;
        RECT 583.930 0.155 592.750 4.280 ;
        RECT 593.590 0.155 602.410 4.280 ;
        RECT 603.250 0.155 612.070 4.280 ;
        RECT 612.910 0.155 621.730 4.280 ;
        RECT 622.570 0.155 631.390 4.280 ;
        RECT 632.230 0.155 641.050 4.280 ;
        RECT 641.890 0.155 650.710 4.280 ;
        RECT 651.550 0.155 660.370 4.280 ;
        RECT 661.210 0.155 670.030 4.280 ;
        RECT 670.870 0.155 679.690 4.280 ;
        RECT 680.530 0.155 689.350 4.280 ;
        RECT 690.190 0.155 699.010 4.280 ;
        RECT 699.850 0.155 708.670 4.280 ;
        RECT 709.510 0.155 718.330 4.280 ;
        RECT 719.170 0.155 727.990 4.280 ;
        RECT 728.830 0.155 737.650 4.280 ;
        RECT 738.490 0.155 747.310 4.280 ;
        RECT 748.150 0.155 756.970 4.280 ;
        RECT 757.810 0.155 766.630 4.280 ;
        RECT 767.470 0.155 776.290 4.280 ;
        RECT 777.130 0.155 785.950 4.280 ;
        RECT 786.790 0.155 799.380 4.280 ;
      LAYER met3 ;
        RECT 1.445 0.175 798.955 636.645 ;
      LAYER met4 ;
        RECT 2.135 10.240 20.640 607.745 ;
        RECT 23.040 10.240 97.440 607.745 ;
        RECT 99.840 10.240 174.240 607.745 ;
        RECT 176.640 10.240 251.040 607.745 ;
        RECT 253.440 10.240 327.840 607.745 ;
        RECT 330.240 10.240 404.640 607.745 ;
        RECT 407.040 10.240 481.440 607.745 ;
        RECT 483.840 10.240 558.240 607.745 ;
        RECT 560.640 10.240 635.040 607.745 ;
        RECT 637.440 10.240 711.840 607.745 ;
        RECT 714.240 10.240 787.225 607.745 ;
        RECT 2.135 2.215 787.225 10.240 ;
  END
END bec
END LIBRARY

