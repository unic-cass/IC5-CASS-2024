magic
tech sky130A
magscale 1 2
timestamp 1731516492
<< nwell >>
rect 1066 106885 108874 107451
rect 1066 105797 108874 106363
rect 1066 104709 108874 105275
rect 1066 103621 108874 104187
rect 1066 102533 108874 103099
rect 1066 101445 108874 102011
rect 1066 100357 108874 100923
rect 1066 99269 108874 99835
rect 1066 98181 108874 98747
rect 1066 97093 108874 97659
rect 1066 96005 108874 96571
rect 1066 94917 108874 95483
rect 1066 93829 108874 94395
rect 1066 92741 108874 93307
rect 1066 91653 108874 92219
rect 1066 90565 108874 91131
rect 1066 89477 108874 90043
rect 1066 88389 108874 88955
rect 1066 87301 108874 87867
rect 1066 86213 108874 86779
rect 1066 85125 108874 85691
rect 1066 84037 108874 84603
rect 1066 82949 108874 83515
rect 1066 81861 108874 82427
rect 1066 80773 108874 81339
rect 1066 79685 108874 80251
rect 1066 78597 108874 79163
rect 1066 77509 108874 78075
rect 1066 76421 108874 76987
rect 1066 75333 108874 75899
rect 1066 74245 108874 74811
rect 1066 73157 108874 73723
rect 1066 72069 108874 72635
rect 1066 70981 108874 71547
rect 1066 69893 108874 70459
rect 1066 68805 108874 69371
rect 1066 67717 108874 68283
rect 1066 66629 108874 67195
rect 1066 65541 108874 66107
rect 1066 64453 108874 65019
rect 1066 63365 108874 63931
rect 1066 62277 108874 62843
rect 1066 61189 108874 61755
rect 1066 60101 108874 60667
rect 1066 59013 108874 59579
rect 1066 57925 108874 58491
rect 1066 56837 108874 57403
rect 1066 55749 108874 56315
rect 1066 54661 108874 55227
rect 1066 53573 108874 54139
rect 1066 52485 108874 53051
rect 1066 51397 108874 51963
rect 1066 50309 108874 50875
rect 1066 49221 108874 49787
rect 1066 48133 108874 48699
rect 1066 47045 108874 47611
rect 1066 45957 108874 46523
rect 1066 44869 108874 45435
rect 1066 43781 108874 44347
rect 1066 42693 108874 43259
rect 1066 41605 108874 42171
rect 1066 40517 108874 41083
rect 1066 39429 108874 39995
rect 1066 38341 108874 38907
rect 1066 37253 108874 37819
rect 1066 36165 108874 36731
rect 1066 35077 108874 35643
rect 1066 33989 108874 34555
rect 1066 32901 108874 33467
rect 1066 31813 108874 32379
rect 1066 30725 108874 31291
rect 1066 29637 108874 30203
rect 1066 28549 108874 29115
rect 1066 27461 108874 28027
rect 1066 26373 108874 26939
rect 1066 25285 108874 25851
rect 1066 24197 108874 24763
rect 1066 23109 108874 23675
rect 1066 22021 108874 22587
rect 1066 20933 108874 21499
rect 1066 19845 108874 20411
rect 1066 18757 108874 19323
rect 1066 17669 108874 18235
rect 1066 16581 108874 17147
rect 1066 15493 108874 16059
rect 1066 14405 108874 14971
rect 1066 13317 108874 13883
rect 1066 12229 108874 12795
rect 1066 11141 108874 11707
rect 1066 10053 108874 10619
rect 1066 8965 108874 9531
rect 1066 7877 108874 8443
rect 1066 6789 108874 7355
rect 1066 5701 108874 6267
rect 1066 4613 108874 5179
rect 1066 3525 108874 4091
rect 1066 2437 108874 3003
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 1104 1436 108896 108112
<< metal2 >>
rect 1122 109200 1178 110000
rect 2502 109200 2558 110000
rect 3882 109200 3938 110000
rect 5262 109200 5318 110000
rect 6642 109200 6698 110000
rect 8022 109200 8078 110000
rect 9402 109200 9458 110000
rect 10782 109200 10838 110000
rect 12162 109200 12218 110000
rect 13542 109200 13598 110000
rect 14922 109200 14978 110000
rect 16302 109200 16358 110000
rect 17682 109200 17738 110000
rect 19062 109200 19118 110000
rect 20442 109200 20498 110000
rect 21822 109200 21878 110000
rect 23202 109200 23258 110000
rect 24582 109200 24638 110000
rect 25962 109200 26018 110000
rect 27342 109200 27398 110000
rect 28722 109200 28778 110000
rect 30102 109200 30158 110000
rect 31482 109200 31538 110000
rect 32862 109200 32918 110000
rect 34242 109200 34298 110000
rect 35622 109200 35678 110000
rect 37002 109200 37058 110000
rect 38382 109200 38438 110000
rect 39762 109200 39818 110000
rect 41142 109200 41198 110000
rect 42522 109200 42578 110000
rect 43902 109200 43958 110000
rect 45282 109200 45338 110000
rect 46662 109200 46718 110000
rect 48042 109200 48098 110000
rect 49422 109200 49478 110000
rect 50802 109200 50858 110000
rect 52182 109200 52238 110000
rect 53562 109200 53618 110000
rect 54942 109200 54998 110000
rect 56322 109200 56378 110000
rect 57702 109200 57758 110000
rect 59082 109200 59138 110000
rect 60462 109200 60518 110000
rect 61842 109200 61898 110000
rect 63222 109200 63278 110000
rect 64602 109200 64658 110000
rect 65982 109200 66038 110000
rect 67362 109200 67418 110000
rect 68742 109200 68798 110000
rect 70122 109200 70178 110000
rect 71502 109200 71558 110000
rect 72882 109200 72938 110000
rect 74262 109200 74318 110000
rect 75642 109200 75698 110000
rect 77022 109200 77078 110000
rect 78402 109200 78458 110000
rect 79782 109200 79838 110000
rect 81162 109200 81218 110000
rect 82542 109200 82598 110000
rect 83922 109200 83978 110000
rect 85302 109200 85358 110000
rect 86682 109200 86738 110000
rect 88062 109200 88118 110000
rect 89442 109200 89498 110000
rect 90822 109200 90878 110000
rect 92202 109200 92258 110000
rect 93582 109200 93638 110000
rect 94962 109200 95018 110000
rect 96342 109200 96398 110000
rect 97722 109200 97778 110000
rect 99102 109200 99158 110000
rect 100482 109200 100538 110000
rect 101862 109200 101918 110000
rect 103242 109200 103298 110000
rect 104622 109200 104678 110000
rect 106002 109200 106058 110000
rect 107382 109200 107438 110000
rect 108762 109200 108818 110000
rect 1122 0 1178 800
rect 2778 0 2834 800
rect 4434 0 4490 800
rect 6090 0 6146 800
rect 7746 0 7802 800
rect 9402 0 9458 800
rect 11058 0 11114 800
rect 12714 0 12770 800
rect 14370 0 14426 800
rect 16026 0 16082 800
rect 17682 0 17738 800
rect 19338 0 19394 800
rect 20994 0 21050 800
rect 22650 0 22706 800
rect 24306 0 24362 800
rect 25962 0 26018 800
rect 27618 0 27674 800
rect 29274 0 29330 800
rect 30930 0 30986 800
rect 32586 0 32642 800
rect 34242 0 34298 800
rect 35898 0 35954 800
rect 37554 0 37610 800
rect 39210 0 39266 800
rect 40866 0 40922 800
rect 42522 0 42578 800
rect 44178 0 44234 800
rect 45834 0 45890 800
rect 47490 0 47546 800
rect 49146 0 49202 800
rect 50802 0 50858 800
rect 52458 0 52514 800
rect 54114 0 54170 800
rect 55770 0 55826 800
rect 57426 0 57482 800
rect 59082 0 59138 800
rect 60738 0 60794 800
rect 62394 0 62450 800
rect 64050 0 64106 800
rect 65706 0 65762 800
rect 67362 0 67418 800
rect 69018 0 69074 800
rect 70674 0 70730 800
rect 72330 0 72386 800
rect 73986 0 74042 800
rect 75642 0 75698 800
rect 77298 0 77354 800
rect 78954 0 79010 800
rect 80610 0 80666 800
rect 82266 0 82322 800
rect 83922 0 83978 800
rect 85578 0 85634 800
rect 87234 0 87290 800
rect 88890 0 88946 800
rect 90546 0 90602 800
rect 92202 0 92258 800
rect 93858 0 93914 800
rect 95514 0 95570 800
rect 97170 0 97226 800
rect 98826 0 98882 800
rect 100482 0 100538 800
rect 102138 0 102194 800
rect 103794 0 103850 800
rect 105450 0 105506 800
rect 107106 0 107162 800
rect 108762 0 108818 800
<< obsm2 >>
rect 1234 109144 2446 109290
rect 2614 109144 3826 109290
rect 3994 109144 5206 109290
rect 5374 109144 6586 109290
rect 6754 109144 7966 109290
rect 8134 109144 9346 109290
rect 9514 109144 10726 109290
rect 10894 109144 12106 109290
rect 12274 109144 13486 109290
rect 13654 109144 14866 109290
rect 15034 109144 16246 109290
rect 16414 109144 17626 109290
rect 17794 109144 19006 109290
rect 19174 109144 20386 109290
rect 20554 109144 21766 109290
rect 21934 109144 23146 109290
rect 23314 109144 24526 109290
rect 24694 109144 25906 109290
rect 26074 109144 27286 109290
rect 27454 109144 28666 109290
rect 28834 109144 30046 109290
rect 30214 109144 31426 109290
rect 31594 109144 32806 109290
rect 32974 109144 34186 109290
rect 34354 109144 35566 109290
rect 35734 109144 36946 109290
rect 37114 109144 38326 109290
rect 38494 109144 39706 109290
rect 39874 109144 41086 109290
rect 41254 109144 42466 109290
rect 42634 109144 43846 109290
rect 44014 109144 45226 109290
rect 45394 109144 46606 109290
rect 46774 109144 47986 109290
rect 48154 109144 49366 109290
rect 49534 109144 50746 109290
rect 50914 109144 52126 109290
rect 52294 109144 53506 109290
rect 53674 109144 54886 109290
rect 55054 109144 56266 109290
rect 56434 109144 57646 109290
rect 57814 109144 59026 109290
rect 59194 109144 60406 109290
rect 60574 109144 61786 109290
rect 61954 109144 63166 109290
rect 63334 109144 64546 109290
rect 64714 109144 65926 109290
rect 66094 109144 67306 109290
rect 67474 109144 68686 109290
rect 68854 109144 70066 109290
rect 70234 109144 71446 109290
rect 71614 109144 72826 109290
rect 72994 109144 74206 109290
rect 74374 109144 75586 109290
rect 75754 109144 76966 109290
rect 77134 109144 78346 109290
rect 78514 109144 79726 109290
rect 79894 109144 81106 109290
rect 81274 109144 82486 109290
rect 82654 109144 83866 109290
rect 84034 109144 85246 109290
rect 85414 109144 86626 109290
rect 86794 109144 88006 109290
rect 88174 109144 89386 109290
rect 89554 109144 90766 109290
rect 90934 109144 92146 109290
rect 92314 109144 93526 109290
rect 93694 109144 94906 109290
rect 95074 109144 96286 109290
rect 96454 109144 97666 109290
rect 97834 109144 99046 109290
rect 99214 109144 100426 109290
rect 100594 109144 101806 109290
rect 101974 109144 103186 109290
rect 103354 109144 104566 109290
rect 104734 109144 105946 109290
rect 106114 109144 107326 109290
rect 107494 109144 108706 109290
rect 1124 856 108816 109144
rect 1234 734 2722 856
rect 2890 734 4378 856
rect 4546 734 6034 856
rect 6202 734 7690 856
rect 7858 734 9346 856
rect 9514 734 11002 856
rect 11170 734 12658 856
rect 12826 734 14314 856
rect 14482 734 15970 856
rect 16138 734 17626 856
rect 17794 734 19282 856
rect 19450 734 20938 856
rect 21106 734 22594 856
rect 22762 734 24250 856
rect 24418 734 25906 856
rect 26074 734 27562 856
rect 27730 734 29218 856
rect 29386 734 30874 856
rect 31042 734 32530 856
rect 32698 734 34186 856
rect 34354 734 35842 856
rect 36010 734 37498 856
rect 37666 734 39154 856
rect 39322 734 40810 856
rect 40978 734 42466 856
rect 42634 734 44122 856
rect 44290 734 45778 856
rect 45946 734 47434 856
rect 47602 734 49090 856
rect 49258 734 50746 856
rect 50914 734 52402 856
rect 52570 734 54058 856
rect 54226 734 55714 856
rect 55882 734 57370 856
rect 57538 734 59026 856
rect 59194 734 60682 856
rect 60850 734 62338 856
rect 62506 734 63994 856
rect 64162 734 65650 856
rect 65818 734 67306 856
rect 67474 734 68962 856
rect 69130 734 70618 856
rect 70786 734 72274 856
rect 72442 734 73930 856
rect 74098 734 75586 856
rect 75754 734 77242 856
rect 77410 734 78898 856
rect 79066 734 80554 856
rect 80722 734 82210 856
rect 82378 734 83866 856
rect 84034 734 85522 856
rect 85690 734 87178 856
rect 87346 734 88834 856
rect 89002 734 90490 856
rect 90658 734 92146 856
rect 92314 734 93802 856
rect 93970 734 95458 856
rect 95626 734 97114 856
rect 97282 734 98770 856
rect 98938 734 100426 856
rect 100594 734 102082 856
rect 102250 734 103738 856
rect 103906 734 105394 856
rect 105562 734 107050 856
rect 107218 734 108706 856
<< metal3 >>
rect 109200 82424 110000 82544
rect 109200 27480 110000 27600
<< obsm3 >>
rect 4061 82624 109200 108085
rect 4061 82344 109120 82624
rect 4061 27680 109200 82344
rect 4061 27400 109120 27680
rect 4061 1667 109200 27400
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 4659 107840 102613 108085
rect 4659 2048 19488 107840
rect 19968 2048 34848 107840
rect 35328 2048 50208 107840
rect 50688 2048 65568 107840
rect 66048 2048 80928 107840
rect 81408 2048 96288 107840
rect 96768 2048 102613 107840
rect 4659 1667 102613 2048
<< labels >>
rlabel metal2 s 14922 109200 14978 110000 6 becStatus[0]
port 1 nsew signal input
rlabel metal2 s 16302 109200 16358 110000 6 becStatus[1]
port 2 nsew signal input
rlabel metal2 s 17682 109200 17738 110000 6 becStatus[2]
port 3 nsew signal input
rlabel metal2 s 19062 109200 19118 110000 6 becStatus[3]
port 4 nsew signal input
rlabel metal2 s 21822 109200 21878 110000 6 data_in[0]
port 5 nsew signal input
rlabel metal2 s 49422 109200 49478 110000 6 data_in[10]
port 6 nsew signal input
rlabel metal2 s 52182 109200 52238 110000 6 data_in[11]
port 7 nsew signal input
rlabel metal2 s 54942 109200 54998 110000 6 data_in[12]
port 8 nsew signal input
rlabel metal2 s 57702 109200 57758 110000 6 data_in[13]
port 9 nsew signal input
rlabel metal2 s 60462 109200 60518 110000 6 data_in[14]
port 10 nsew signal input
rlabel metal2 s 63222 109200 63278 110000 6 data_in[15]
port 11 nsew signal input
rlabel metal2 s 65982 109200 66038 110000 6 data_in[16]
port 12 nsew signal input
rlabel metal2 s 68742 109200 68798 110000 6 data_in[17]
port 13 nsew signal input
rlabel metal2 s 71502 109200 71558 110000 6 data_in[18]
port 14 nsew signal input
rlabel metal2 s 74262 109200 74318 110000 6 data_in[19]
port 15 nsew signal input
rlabel metal2 s 24582 109200 24638 110000 6 data_in[1]
port 16 nsew signal input
rlabel metal2 s 77022 109200 77078 110000 6 data_in[20]
port 17 nsew signal input
rlabel metal2 s 79782 109200 79838 110000 6 data_in[21]
port 18 nsew signal input
rlabel metal2 s 82542 109200 82598 110000 6 data_in[22]
port 19 nsew signal input
rlabel metal2 s 85302 109200 85358 110000 6 data_in[23]
port 20 nsew signal input
rlabel metal2 s 88062 109200 88118 110000 6 data_in[24]
port 21 nsew signal input
rlabel metal2 s 90822 109200 90878 110000 6 data_in[25]
port 22 nsew signal input
rlabel metal2 s 93582 109200 93638 110000 6 data_in[26]
port 23 nsew signal input
rlabel metal2 s 96342 109200 96398 110000 6 data_in[27]
port 24 nsew signal input
rlabel metal2 s 99102 109200 99158 110000 6 data_in[28]
port 25 nsew signal input
rlabel metal2 s 101862 109200 101918 110000 6 data_in[29]
port 26 nsew signal input
rlabel metal2 s 27342 109200 27398 110000 6 data_in[2]
port 27 nsew signal input
rlabel metal2 s 104622 109200 104678 110000 6 data_in[30]
port 28 nsew signal input
rlabel metal2 s 107382 109200 107438 110000 6 data_in[31]
port 29 nsew signal input
rlabel metal2 s 30102 109200 30158 110000 6 data_in[3]
port 30 nsew signal input
rlabel metal2 s 32862 109200 32918 110000 6 data_in[4]
port 31 nsew signal input
rlabel metal2 s 35622 109200 35678 110000 6 data_in[5]
port 32 nsew signal input
rlabel metal2 s 38382 109200 38438 110000 6 data_in[6]
port 33 nsew signal input
rlabel metal2 s 41142 109200 41198 110000 6 data_in[7]
port 34 nsew signal input
rlabel metal2 s 43902 109200 43958 110000 6 data_in[8]
port 35 nsew signal input
rlabel metal2 s 46662 109200 46718 110000 6 data_in[9]
port 36 nsew signal input
rlabel metal2 s 23202 109200 23258 110000 6 data_out[0]
port 37 nsew signal output
rlabel metal2 s 50802 109200 50858 110000 6 data_out[10]
port 38 nsew signal output
rlabel metal2 s 53562 109200 53618 110000 6 data_out[11]
port 39 nsew signal output
rlabel metal2 s 56322 109200 56378 110000 6 data_out[12]
port 40 nsew signal output
rlabel metal2 s 59082 109200 59138 110000 6 data_out[13]
port 41 nsew signal output
rlabel metal2 s 61842 109200 61898 110000 6 data_out[14]
port 42 nsew signal output
rlabel metal2 s 64602 109200 64658 110000 6 data_out[15]
port 43 nsew signal output
rlabel metal2 s 67362 109200 67418 110000 6 data_out[16]
port 44 nsew signal output
rlabel metal2 s 70122 109200 70178 110000 6 data_out[17]
port 45 nsew signal output
rlabel metal2 s 72882 109200 72938 110000 6 data_out[18]
port 46 nsew signal output
rlabel metal2 s 75642 109200 75698 110000 6 data_out[19]
port 47 nsew signal output
rlabel metal2 s 25962 109200 26018 110000 6 data_out[1]
port 48 nsew signal output
rlabel metal2 s 78402 109200 78458 110000 6 data_out[20]
port 49 nsew signal output
rlabel metal2 s 81162 109200 81218 110000 6 data_out[21]
port 50 nsew signal output
rlabel metal2 s 83922 109200 83978 110000 6 data_out[22]
port 51 nsew signal output
rlabel metal2 s 86682 109200 86738 110000 6 data_out[23]
port 52 nsew signal output
rlabel metal2 s 89442 109200 89498 110000 6 data_out[24]
port 53 nsew signal output
rlabel metal2 s 92202 109200 92258 110000 6 data_out[25]
port 54 nsew signal output
rlabel metal2 s 94962 109200 95018 110000 6 data_out[26]
port 55 nsew signal output
rlabel metal2 s 97722 109200 97778 110000 6 data_out[27]
port 56 nsew signal output
rlabel metal2 s 100482 109200 100538 110000 6 data_out[28]
port 57 nsew signal output
rlabel metal2 s 103242 109200 103298 110000 6 data_out[29]
port 58 nsew signal output
rlabel metal2 s 28722 109200 28778 110000 6 data_out[2]
port 59 nsew signal output
rlabel metal2 s 106002 109200 106058 110000 6 data_out[30]
port 60 nsew signal output
rlabel metal2 s 108762 109200 108818 110000 6 data_out[31]
port 61 nsew signal output
rlabel metal2 s 31482 109200 31538 110000 6 data_out[3]
port 62 nsew signal output
rlabel metal2 s 34242 109200 34298 110000 6 data_out[4]
port 63 nsew signal output
rlabel metal2 s 37002 109200 37058 110000 6 data_out[5]
port 64 nsew signal output
rlabel metal2 s 39762 109200 39818 110000 6 data_out[6]
port 65 nsew signal output
rlabel metal2 s 42522 109200 42578 110000 6 data_out[7]
port 66 nsew signal output
rlabel metal2 s 45282 109200 45338 110000 6 data_out[8]
port 67 nsew signal output
rlabel metal2 s 48042 109200 48098 110000 6 data_out[9]
port 68 nsew signal output
rlabel metal3 s 109200 82424 110000 82544 6 io_oeb
port 69 nsew signal output
rlabel metal3 s 109200 27480 110000 27600 6 io_out
port 70 nsew signal output
rlabel metal2 s 10782 109200 10838 110000 6 ki
port 71 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 la_data_in[0]
port 72 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[10]
port 73 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[11]
port 74 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[12]
port 75 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[13]
port 76 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[14]
port 77 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[15]
port 78 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[16]
port 79 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[17]
port 80 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[18]
port 81 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[19]
port 82 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la_data_in[1]
port 83 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[20]
port 84 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[21]
port 85 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[22]
port 86 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[23]
port 87 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[24]
port 88 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[25]
port 89 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[26]
port 90 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[27]
port 91 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[28]
port 92 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_data_in[29]
port 93 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 la_data_in[2]
port 94 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[30]
port 95 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[31]
port 96 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 la_data_in[3]
port 97 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 la_data_in[4]
port 98 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 la_data_in[5]
port 99 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[6]
port 100 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[7]
port 101 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[8]
port 102 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[9]
port 103 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 la_data_out[0]
port 104 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[10]
port 105 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[11]
port 106 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[12]
port 107 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[13]
port 108 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[14]
port 109 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[15]
port 110 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[16]
port 111 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[17]
port 112 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[18]
port 113 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[19]
port 114 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 la_data_out[1]
port 115 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[20]
port 116 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[21]
port 117 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[22]
port 118 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[23]
port 119 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[24]
port 120 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[25]
port 121 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[26]
port 122 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[27]
port 123 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[28]
port 124 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[29]
port 125 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 la_data_out[2]
port 126 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[30]
port 127 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[31]
port 128 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 la_data_out[3]
port 129 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[4]
port 130 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 la_data_out[5]
port 131 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[6]
port 132 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 la_data_out[7]
port 133 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[8]
port 134 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 la_data_out[9]
port 135 nsew signal output
rlabel metal2 s 9402 109200 9458 110000 6 load_data
port 136 nsew signal output
rlabel metal2 s 1122 109200 1178 110000 6 load_status[0]
port 137 nsew signal output
rlabel metal2 s 2502 109200 2558 110000 6 load_status[1]
port 138 nsew signal output
rlabel metal2 s 3882 109200 3938 110000 6 load_status[2]
port 139 nsew signal output
rlabel metal2 s 5262 109200 5318 110000 6 load_status[3]
port 140 nsew signal output
rlabel metal2 s 6642 109200 6698 110000 6 load_status[4]
port 141 nsew signal output
rlabel metal2 s 8022 109200 8078 110000 6 load_status[5]
port 142 nsew signal output
rlabel metal2 s 12162 109200 12218 110000 6 next_key
port 143 nsew signal input
rlabel metal2 s 13542 109200 13598 110000 6 slv_done
port 144 nsew signal input
rlabel metal2 s 20442 109200 20498 110000 6 slv_enable
port 145 nsew signal output
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 146 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 147 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 147 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 147 nsew ground bidirectional
rlabel metal2 s 1122 0 1178 800 6 wb_clk_i
port 148 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wb_rst_i
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38506586
string GDS_FILE /home/cass/projects/IC5-CASS-2024/openlane/lovers_controller/runs/24_11_13_23_23/results/signoff/lovers_controller.magic.gds
string GDS_START 625646
<< end >>

