* NGSPICE file created from vmsu_8bit_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt vmsu_8bit_top a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] b[0] b[1] b[2] b[3]
+ b[4] b[5] b[6] b[7] clk control p[0] p[10] p[11] p[12] p[13] p[14] p[15] p[1] p[2]
+ p[3] p[4] p[5] p[6] p[7] p[8] p[9] rst vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1605__44 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1676_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_40_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1620__58 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1690_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1270_ _1274_/A _1273_/B _1259_/X _1267_/Y vssd1 vssd1 vccd1 vccd1 _1270_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0985_ _0985_/A _0985_/B vssd1 vssd1 vccd1 vccd1 _0986_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1468_ hold98/X vssd1 vssd1 vccd1 vccd1 _1694_/D sky130_fd_sc_hd__clkbuf_1
X_1399_ _1399_/A vssd1 vssd1 vccd1 vccd1 _1709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1537_ _1537_/A hold41/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1596__35 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1667_/CLK sky130_fd_sc_hd__inv_2
X_1253_ _1245_/B _1249_/A _1244_/B vssd1 vssd1 vccd1 vccd1 _1288_/C sky130_fd_sc_hd__o21a_1
X_1322_ _1327_/A _1323_/B _1323_/A vssd1 vssd1 vccd1 vccd1 _1324_/A sky130_fd_sc_hd__nand3_1
X_1184_ _1220_/B _1221_/A _1221_/B vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0968_ _1106_/A _1107_/A vssd1 vssd1 vccd1 vccd1 _1062_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0899_ _0899_/A _0899_/B vssd1 vssd1 vccd1 vccd1 _0900_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1305_ _1330_/B _1305_/B vssd1 vssd1 vccd1 vccd1 _1314_/B sky130_fd_sc_hd__and2_1
X_1236_ _1236_/A _1236_/B vssd1 vssd1 vccd1 vccd1 _1361_/B sky130_fd_sc_hd__nor2_1
X_1167_ _1167_/A vssd1 vssd1 vccd1 vccd1 _1168_/C sky130_fd_sc_hd__inv_2
X_1098_ _1098_/A _1098_/B _1098_/C vssd1 vssd1 vccd1 vccd1 _1103_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1021_ _1021_/A vssd1 vssd1 vccd1 vccd1 _1022_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1219_ _1364_/C _1219_/B vssd1 vssd1 vccd1 vccd1 _1236_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_1626__64 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1696_/CLK sky130_fd_sc_hd__inv_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__inv_2
XFILLER_0_44_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1004_ _1345_/B _1004_/B vssd1 vssd1 vccd1 vccd1 _1347_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1699_ _1699_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _1699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput20 _1695_/Q vssd1 vssd1 vccd1 vccd1 p[10] sky130_fd_sc_hd__buf_12
Xoutput31 _1691_/Q vssd1 vssd1 vccd1 vccd1 p[6] sky130_fd_sc_hd__buf_12
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ hold13/X hold2/X _1577_/A vssd1 vssd1 vccd1 vccd1 _1553_/X sky130_fd_sc_hd__or3_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ _1482_/Y hold28/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__a21oi_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0984_ _0984_/A vssd1 vssd1 vccd1 vccd1 _1347_/A sky130_fd_sc_hd__inv_2
X_1536_ hold41/X _1537_/A vssd1 vssd1 vccd1 vccd1 _1538_/A sky130_fd_sc_hd__or2_1
X_1398_ _1588_/B input8/X vssd1 vssd1 vccd1 vccd1 _1399_/A sky130_fd_sc_hd__and2_1
X_1467_ _1467_/A _1588_/B hold97/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__and3_1
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1252_ _1290_/A _1252_/B _1252_/C vssd1 vssd1 vccd1 vccd1 _1295_/C sky130_fd_sc_hd__nand3_2
X_1321_ _1321_/A _1330_/C vssd1 vssd1 vccd1 vccd1 _1323_/B sky130_fd_sc_hd__nand2_1
X_1183_ _1209_/B _1208_/A _1208_/B vssd1 vssd1 vccd1 vccd1 _1221_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0967_ _1682_/Q _1668_/Q vssd1 vssd1 vccd1 vccd1 _1107_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1519_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1680_/D sky130_fd_sc_hd__clkbuf_1
X_0898_ _0898_/A vssd1 vssd1 vccd1 vccd1 _0909_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1166_ _1166_/A _1167_/A vssd1 vssd1 vccd1 vccd1 _1172_/A sky130_fd_sc_hd__nand2_1
X_1235_ _1414_/A _1231_/Y _1234_/Y vssd1 vssd1 vccd1 vccd1 _1236_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1304_ _1667_/Q _1676_/Q _1668_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1305_/B sky130_fd_sc_hd__a22o_1
X_1097_ _1097_/A _1097_/B vssd1 vssd1 vccd1 vccd1 _1158_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ _1020_/A vssd1 vssd1 vccd1 vccd1 _1022_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1149_ _1149_/A _1149_/B vssd1 vssd1 vccd1 vccd1 _1151_/A sky130_fd_sc_hd__nand2_1
X_1218_ _1218_/A _1218_/B vssd1 vssd1 vccd1 vccd1 _1219_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1654__4 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1724_/CLK sky130_fd_sc_hd__inv_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1641__24 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1711_/CLK sky130_fd_sc_hd__inv_2
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1003_ _1003_/A _1004_/B _1003_/C vssd1 vssd1 vccd1 vccd1 _1345_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_44_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1698_ _1698_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 _1698_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput21 _1696_/Q vssd1 vssd1 vccd1 vccd1 p[11] sky130_fd_sc_hd__buf_12
Xoutput32 _1692_/Q vssd1 vssd1 vccd1 vccd1 p[7] sky130_fd_sc_hd__buf_12
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1552_ _1592_/A hold2/X vssd1 vssd1 vccd1 vccd1 _1674_/D sky130_fd_sc_hd__nor2_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _1506_/A hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__nand2_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _0983_/A _1351_/B vssd1 vssd1 vccd1 vccd1 _0984_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1535_ hold37/A _1541_/B vssd1 vssd1 vccd1 vccd1 _1537_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1397_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1710_/D sky130_fd_sc_hd__clkbuf_1
X_1466_ hold88/X hold16/X hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__a21o_1
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ _1320_/A _1320_/B vssd1 vssd1 vccd1 vccd1 _1330_/C sky130_fd_sc_hd__nand2_1
X_1182_ _1182_/A _1182_/B vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__nand2_1
X_1251_ _1251_/A _1251_/B vssd1 vssd1 vccd1 vccd1 _1252_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0966_ _1680_/Q _1670_/Q vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__nand2_1
X_0897_ _0899_/A _0899_/B vssd1 vssd1 vccd1 vccd1 _0898_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1449_ _1506_/A hold24/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__nand2_1
X_1518_ _1518_/A _1588_/B hold65/X vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__and3_1
XFILLER_0_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1303_ _1303_/A _1303_/B _1303_/C _1303_/D vssd1 vssd1 vccd1 vccd1 _1330_/B sky130_fd_sc_hd__or4_1
XFILLER_0_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1165_ _1239_/B _1165_/B vssd1 vssd1 vccd1 vccd1 _1167_/A sky130_fd_sc_hd__nand2_1
X_1096_ _1098_/B vssd1 vssd1 vccd1 vccd1 _1097_/B sky130_fd_sc_hd__inv_2
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1234_ _1414_/B vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__inv_2
X_1647__30 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1717_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0949_ _0953_/A _0953_/B vssd1 vssd1 vccd1 vccd1 _0989_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1148_ _1148_/A _1200_/A _1148_/C vssd1 vssd1 vccd1 vccd1 _1199_/A sky130_fd_sc_hd__nand3_1
X_1079_ _1079_/A _1079_/B _1079_/C vssd1 vssd1 vccd1 vccd1 _1083_/A sky130_fd_sc_hd__nand3_1
X_1217_ _1301_/B vssd1 vssd1 vccd1 vccd1 _1364_/C sky130_fd_sc_hd__inv_2
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1002_ _1342_/C vssd1 vssd1 vccd1 vccd1 _1003_/C sky130_fd_sc_hd__inv_2
XFILLER_0_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1617__55 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1687_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1697_ _1697_/CLK hold23/X vssd1 vssd1 vccd1 vccd1 _1697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput33 _1693_/Q vssd1 vssd1 vccd1 vccd1 p[8] sky130_fd_sc_hd__buf_12
Xoutput22 _1697_/Q vssd1 vssd1 vccd1 vccd1 p[12] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1551_ hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__inv_2
X_1482_ _1425_/B _1425_/A _1479_/A vssd1 vssd1 vccd1 vccd1 _1482_/Y sky130_fd_sc_hd__o21ai_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0982_ _0982_/A _0982_/B _0982_/C vssd1 vssd1 vccd1 vccd1 _1351_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1465_ hold17/A _1506_/A hold96/X vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__or3b_1
X_1534_ hold44/X _1534_/B vssd1 vssd1 vccd1 vccd1 _1541_/B sky130_fd_sc_hd__nor2_1
X_1396_ _1588_/B input9/X vssd1 vssd1 vccd1 vccd1 _1397_/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1250_ _1250_/A _1250_/B vssd1 vssd1 vccd1 vccd1 _1290_/A sky130_fd_sc_hd__nand2_1
X_1181_ _1208_/B vssd1 vssd1 vccd1 vccd1 _1182_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0965_ _1036_/C _0965_/B vssd1 vssd1 vccd1 vccd1 _0977_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0896_ _0896_/A _1681_/Q _1671_/Q vssd1 vssd1 vccd1 vccd1 _0899_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1448_ hold88/X vssd1 vssd1 vccd1 vccd1 _1506_/A sky130_fd_sc_hd__inv_2
X_1517_ hold37/A _1521_/A hold64/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__o21ai_1
X_1379_ _1592_/A _1577_/A vssd1 vssd1 vccd1 vccd1 _1719_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_45_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1233_ _1233_/A _1233_/B _1233_/C vssd1 vssd1 vccd1 vccd1 _1414_/B sky130_fd_sc_hd__nand3_1
X_1302_ _1302_/A _1302_/B _1302_/C vssd1 vssd1 vccd1 vccd1 _1376_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_19_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1095_ _1156_/A _1095_/B vssd1 vssd1 vccd1 vccd1 _1098_/B sky130_fd_sc_hd__nand2_1
X_1164_ _1671_/Q _1676_/Q _1672_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1165_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_35_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0948_ _1064_/B _0948_/B vssd1 vssd1 vccd1 vccd1 _0953_/B sky130_fd_sc_hd__nand2_1
X_1662__12 _1613_/A vssd1 vssd1 vccd1 vccd1 _1732_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0879_ _0902_/A _0879_/B _0879_/C vssd1 vssd1 vccd1 vccd1 _0901_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1216_ _1218_/B _1218_/A vssd1 vssd1 vccd1 vccd1 _1301_/B sky130_fd_sc_hd__nor2_1
X_1147_ _1151_/B vssd1 vssd1 vccd1 vccd1 _1148_/C sky130_fd_sc_hd__inv_2
X_1078_ _1078_/A _1078_/B vssd1 vssd1 vccd1 vccd1 _1080_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1001_ _1341_/B _1341_/A vssd1 vssd1 vccd1 vccd1 _1342_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1696_ _1696_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 _1696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput34 _1683_/Q vssd1 vssd1 vccd1 vccd1 p[9] sky130_fd_sc_hd__buf_12
Xoutput23 _1698_/Q vssd1 vssd1 vccd1 vccd1 p[13] sky130_fd_sc_hd__buf_12
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1481_ hold91/X vssd1 vssd1 vccd1 vccd1 _1691_/D sky130_fd_sc_hd__clkbuf_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _1548_/Y _1549_/Y _1588_/B hold8/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__o211a_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1679_ _1679_/CLK _1679_/D vssd1 vssd1 vccd1 vccd1 _1679_/Q sky130_fd_sc_hd__dfxtp_4
X_0981_ _0981_/A vssd1 vssd1 vccd1 vccd1 _0982_/C sky130_fd_sc_hd__inv_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0138_ clkbuf_0__0138_/X vssd1 vssd1 vccd1 vccd1 _1644__27/A sky130_fd_sc_hd__clkbuf_16
X_1395_ _1395_/A vssd1 vssd1 vccd1 vccd1 _1711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1464_ hold16/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__inv_2
X_1533_ hold46/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1601__40 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1672_/CLK sky130_fd_sc_hd__inv_2
X_1180_ _1180_/A _1180_/B vssd1 vssd1 vccd1 vccd1 _1208_/B sky130_fd_sc_hd__nand2_1
X_0964_ _0964_/A _0964_/B vssd1 vssd1 vccd1 vccd1 _0965_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1516_ hold64/X hold37/A _1521_/A vssd1 vssd1 vccd1 vccd1 _1518_/A sky130_fd_sc_hd__or3_1
X_0895_ _0895_/A _1679_/Q _1673_/Q vssd1 vssd1 vccd1 vccd1 _0899_/A sky130_fd_sc_hd__nand3_1
X_1378_ hold36/A hold3/X vssd1 vssd1 vccd1 vccd1 _1577_/A sky130_fd_sc_hd__nand2_2
X_1447_ hold24/X _1437_/B _1445_/A vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1232_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1233_/C sky130_fd_sc_hd__inv_2
X_1301_ _1301_/A _1301_/B vssd1 vssd1 vccd1 vccd1 _1302_/C sky130_fd_sc_hd__nand2_1
X_1094_ _1159_/C _1094_/B _1094_/C vssd1 vssd1 vccd1 vccd1 _1095_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1163_ _1163_/A _1163_/B _1303_/C _1303_/D vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__or4_2
X_0947_ _0945_/A _1260_/A _0945_/C vssd1 vssd1 vccd1 vccd1 _0948_/B sky130_fd_sc_hd__o21ai_1
X_0878_ _0911_/C _0888_/A vssd1 vssd1 vccd1 vccd1 _0886_/A sky130_fd_sc_hd__nand2_1
X_1638__21 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1708_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1146_ _1150_/A _1197_/A _1149_/B vssd1 vssd1 vccd1 vccd1 _1200_/A sky130_fd_sc_hd__nand3_1
X_1215_ _1215_/A _1291_/B vssd1 vssd1 vccd1 vccd1 _1218_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1077_ _1079_/A vssd1 vssd1 vccd1 vccd1 _1078_/B sky130_fd_sc_hd__inv_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1000_ _1000_/A _1000_/B vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1695_ _1695_/CLK _1695_/D vssd1 vssd1 vccd1 vccd1 _1695_/Q sky130_fd_sc_hd__dfxtp_1
X_1129_ _1129_/A _1129_/B vssd1 vssd1 vccd1 vccd1 _1229_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput24 _1699_/Q vssd1 vssd1 vccd1 vccd1 p[14] sky130_fd_sc_hd__buf_12
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1622__60 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1692_/CLK sky130_fd_sc_hd__inv_2
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1480_/A _1588_/B hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__and3_1
XFILLER_0_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1678_ _1678_/CLK hold47/X vssd1 vssd1 vccd1 vccd1 _1678_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ _0980_/A _0981_/A vssd1 vssd1 vccd1 vccd1 _0983_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1532_ hold45/X _1588_/B _1532_/C vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__and3_1
XFILLER_0_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1463_ hold79/X vssd1 vssd1 vccd1 vccd1 _1695_/D sky130_fd_sc_hd__clkbuf_1
X_1394_ _1588_/B _1394_/B vssd1 vssd1 vccd1 vccd1 _1395_/A sky130_fd_sc_hd__and2_1
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ _0964_/B _0964_/A vssd1 vssd1 vccd1 vccd1 _1036_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_24_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0894_ _1339_/B _1337_/B vssd1 vssd1 vccd1 vccd1 _0905_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1515_ _1702_/Q hold10/X vssd1 vssd1 vccd1 vccd1 _1521_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1446_ _1444_/X hold6/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__a21oi_1
X_1377_ _1375_/Y _1376_/Y _1592_/A vssd1 vssd1 vccd1 vccd1 _1720_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1657__7 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1727_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1231_ _1416_/B vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__inv_2
X_1162_ _1675_/Q vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__inv_2
X_1300_ _1370_/C _1299_/Y _1289_/A vssd1 vssd1 vccd1 vccd1 _1302_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ _1094_/B _1159_/C vssd1 vssd1 vccd1 vccd1 _1156_/A sky130_fd_sc_hd__or2_1
XFILLER_0_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0946_ _0946_/A vssd1 vssd1 vccd1 vccd1 _1064_/B sky130_fd_sc_hd__inv_2
X_0877_ _0879_/C vssd1 vssd1 vccd1 vccd1 _0888_/A sky130_fd_sc_hd__inv_2
XFILLER_0_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1429_ hold18/X hold82/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1145_ _1150_/C vssd1 vssd1 vccd1 vccd1 _1149_/B sky130_fd_sc_hd__inv_2
X_1214_ _1214_/A _1252_/B _1214_/C vssd1 vssd1 vccd1 vccd1 _1291_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_1_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1076_ _1076_/A _1076_/B vssd1 vssd1 vccd1 vccd1 _1079_/A sky130_fd_sc_hd__nand2_1
X_0929_ _0929_/A _1679_/Q _1671_/Q vssd1 vssd1 vccd1 vccd1 _0932_/B sky130_fd_sc_hd__and3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__buf_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1694_ _1694_/CLK _1694_/D vssd1 vssd1 vccd1 vccd1 _1694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1059_ _1059_/A _1059_/B vssd1 vssd1 vccd1 vccd1 _1062_/B sky130_fd_sc_hd__nand2_1
X_1128_ _1128_/A _1178_/A vssd1 vssd1 vccd1 vccd1 _1129_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1608__47 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1679_/CLK sky130_fd_sc_hd__inv_2
Xoutput25 _1686_/Q vssd1 vssd1 vccd1 vccd1 p[15] sky130_fd_sc_hd__buf_12
XFILLER_0_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1677_ _1677_/CLK _1677_/D vssd1 vssd1 vccd1 vccd1 _1677_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1599__38 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1670_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1462_ _1462_/A _1588_/B hold78/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__and3_1
X_1531_ _1534_/B hold44/X _1543_/B vssd1 vssd1 vccd1 vccd1 _1532_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1393_ _1393_/A vssd1 vssd1 vccd1 vccd1 _1712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1729_ _1729_/CLK _1729_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0962_ _1263_/D _0962_/B _0999_/A vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0893_ _1337_/A _1337_/B _1333_/A vssd1 vssd1 vccd1 vccd1 _1339_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1514_ hold63/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__inv_2
X_1445_ _1445_/A hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1376_ _1376_/A _1376_/B _1376_/C vssd1 vssd1 vccd1 vccd1 _1376_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1092_ _1092_/A _1156_/B vssd1 vssd1 vccd1 vccd1 _1159_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1230_ _1230_/A _1230_/B _1230_/C vssd1 vssd1 vccd1 vccd1 _1416_/B sky130_fd_sc_hd__nand3_2
X_1161_ _1676_/Q vssd1 vssd1 vccd1 vccd1 _1303_/C sky130_fd_sc_hd__inv_2
XFILLER_0_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0945_ _0945_/A _1260_/A _0945_/C vssd1 vssd1 vccd1 vccd1 _0946_/A sky130_fd_sc_hd__nor3_1
X_0876_ _0895_/A _0896_/A vssd1 vssd1 vccd1 vccd1 _0879_/C sky130_fd_sc_hd__nor2_1
X_1428_ hold81/X hold49/A vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__nand2_1
X_1359_ _1359_/A _1588_/B _1359_/C vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__and3_1
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1629__67 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1699_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1213_ _1251_/B vssd1 vssd1 vccd1 vccd1 _1214_/A sky130_fd_sc_hd__inv_2
X_1144_ _1149_/A _1150_/C vssd1 vssd1 vccd1 vccd1 _1148_/A sky130_fd_sc_hd__nand2_1
X_1075_ _1071_/A _1074_/Y _1073_/B vssd1 vssd1 vccd1 vccd1 _1076_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0859_ _0868_/A _0869_/A vssd1 vssd1 vccd1 vccd1 _0907_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ _0985_/A _0985_/B _0928_/C vssd1 vssd1 vccd1 vccd1 _0995_/B sky130_fd_sc_hd__nand3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1693_ _1693_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _1693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ _1131_/B _1058_/B vssd1 vssd1 vccd1 vccd1 _1059_/B sky130_fd_sc_hd__nand2_1
X_1127_ _1178_/A _1128_/A vssd1 vssd1 vccd1 vccd1 _1129_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput26 _1694_/Q vssd1 vssd1 vccd1 vccd1 p[1] sky130_fd_sc_hd__buf_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1676_ _1676_/CLK _1676_/D vssd1 vssd1 vccd1 vccd1 _1676_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1392_ _1588_/B _1392_/B vssd1 vssd1 vccd1 vccd1 _1393_/A sky130_fd_sc_hd__and2_1
X_1461_ _1461_/A hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__nand2_1
X_1530_ _1534_/B _1543_/B hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__a21o_1
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold100 _1421_/B vssd1 vssd1 vccd1 vccd1 _1492_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _1728_/CLK _1728_/D vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0961_ _1030_/B _0961_/B vssd1 vssd1 vccd1 vccd1 _0964_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0892_ _1334_/B _1334_/A vssd1 vssd1 vccd1 vccd1 _1333_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1444_ hold5/X _1445_/A vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__or2_1
X_1513_ _1511_/X hold11/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__a21oi_1
X_1375_ _1375_/A _1375_/B vssd1 vssd1 vccd1 vccd1 _1375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1160_ _1168_/A _1188_/A vssd1 vssd1 vccd1 vccd1 _1166_/A sky130_fd_sc_hd__nand2_1
X_1091_ _1091_/A _1091_/B vssd1 vssd1 vccd1 vccd1 _1156_/B sky130_fd_sc_hd__nand2_1
X_0944_ _1681_/Q _1670_/Q vssd1 vssd1 vccd1 vccd1 _0945_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0875_ _1682_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _0896_/A sky130_fd_sc_hd__nand2_1
X_1427_ hold48/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__inv_2
X_1358_ _1358_/A _1358_/B vssd1 vssd1 vccd1 vccd1 _1359_/C sky130_fd_sc_hd__nand2_1
X_1289_ _1289_/A _1299_/A vssd1 vssd1 vccd1 vccd1 _1369_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1644__27 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1714_/CLK sky130_fd_sc_hd__inv_2
X_1212_ _1233_/B _1251_/B vssd1 vssd1 vccd1 vccd1 _1215_/A sky130_fd_sc_hd__nand2_1
X_1143_ _1241_/B _1143_/B vssd1 vssd1 vccd1 vccd1 _1150_/C sky130_fd_sc_hd__nand2_1
X_1074_ _1074_/A vssd1 vssd1 vccd1 vccd1 _1074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0927_ _0997_/B vssd1 vssd1 vccd1 vccd1 _0928_/C sky130_fd_sc_hd__inv_2
X_0858_ _1682_/Q _1671_/Q vssd1 vssd1 vccd1 vccd1 _0869_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1692_ _1692_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 _1692_/Q sky130_fd_sc_hd__dfxtp_1
X_1126_ _1179_/A _1126_/B vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__nor2_1
X_1057_ _1057_/A _1057_/B vssd1 vssd1 vccd1 vccd1 _1131_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput27 _1687_/Q vssd1 vssd1 vccd1 vccd1 p[2] sky130_fd_sc_hd__buf_12
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1675_ _1675_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _1675_/Q sky130_fd_sc_hd__dfxtp_2
X_1109_ _1109_/A _1109_/B vssd1 vssd1 vccd1 vccd1 _1134_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1391_ _1391_/A vssd1 vssd1 vccd1 vccd1 _1713_/D sky130_fd_sc_hd__clkbuf_1
X_1460_ hold77/X _1461_/A vssd1 vssd1 vccd1 vccd1 _1462_/A sky130_fd_sc_hd__or2_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold101 _1702_/Q vssd1 vssd1 vccd1 vccd1 _1508_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1727_ _1727_/CLK _1727_/D vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1589_ hold76/X vssd1 vssd1 vccd1 vccd1 _1668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ _1088_/A _1089_/A vssd1 vssd1 vccd1 vccd1 _0961_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0891_ _0972_/A _0962_/B _0891_/C vssd1 vssd1 vccd1 vccd1 _1334_/A sky130_fd_sc_hd__or3_1
X_1512_ _1511_/B hold37/A hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1443_ _1496_/B hold88/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__nand2_1
X_1374_ _1700_/Q _1374_/B _1375_/A vssd1 vssd1 vccd1 vccd1 _1721_/D sky130_fd_sc_hd__nor3b_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1090_ _1091_/A _1091_/B vssd1 vssd1 vccd1 vccd1 _1092_/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0943_ _1682_/Q vssd1 vssd1 vccd1 vccd1 _0945_/A sky130_fd_sc_hd__inv_2
X_0874_ _1680_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _0895_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1288_ _1295_/C _1288_/B _1288_/C vssd1 vssd1 vccd1 vccd1 _1299_/A sky130_fd_sc_hd__nand3_1
X_1426_ hold80/X _1476_/A vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__nor2_1
X_1357_ _1357_/A vssd1 vssd1 vccd1 vccd1 _1726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1211_ _1211_/A _1211_/B vssd1 vssd1 vccd1 vccd1 _1251_/B sky130_fd_sc_hd__nand2_1
X_1142_ _1667_/Q _1680_/Q _1668_/Q _1679_/Q vssd1 vssd1 vccd1 vccd1 _1143_/B sky130_fd_sc_hd__a22o_1
X_1073_ _1073_/A _1073_/B vssd1 vssd1 vccd1 vccd1 _1076_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0857_ _1681_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _0868_/A sky130_fd_sc_hd__nand2_1
X_0926_ _0926_/A _0926_/B _0926_/C vssd1 vssd1 vccd1 vccd1 _0997_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1704_/D sky130_fd_sc_hd__clkbuf_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__buf_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1691_ _1691_/CLK _1691_/D vssd1 vssd1 vccd1 vccd1 _1691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1125_ _1178_/B vssd1 vssd1 vccd1 vccd1 _1126_/B sky130_fd_sc_hd__inv_2
X_1056_ _1056_/A vssd1 vssd1 vccd1 vccd1 _1057_/B sky130_fd_sc_hd__inv_2
XFILLER_0_35_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0909_ _0909_/A _0909_/B _0911_/A vssd1 vssd1 vccd1 vccd1 _0910_/B sky130_fd_sc_hd__and3_1
Xoutput28 _1688_/Q vssd1 vssd1 vccd1 vccd1 p[3] sky130_fd_sc_hd__buf_12
XFILLER_0_22_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1674_ _1674_/CLK _1674_/D vssd1 vssd1 vccd1 vccd1 _1674_/Q sky130_fd_sc_hd__dfxtp_2
X_1108_ _1109_/A _1109_/B vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__or2_1
X_1039_ _1679_/Q _1670_/Q vssd1 vssd1 vccd1 vccd1 _1052_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1390_ _1588_/B _1390_/B vssd1 vssd1 vccd1 vccd1 _1391_/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 _1719_/Q vssd1 vssd1 vccd1 vccd1 _0834_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _1588_/A _1588_/B hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__and3_1
X_1726_ _1726_/CLK _1726_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0890_ _1673_/Q vssd1 vssd1 vccd1 vccd1 _0962_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1442_ _1442_/A hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__nand2_2
X_1511_ hold10/X _1511_/B hold37/A vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1373_ _1376_/A _1376_/B vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__nand2_1
X_1665__15 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1735_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1709_ _1709_/CLK _1709_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0942_ _1033_/B _0942_/B vssd1 vssd1 vccd1 vccd1 _0953_/A sky130_fd_sc_hd__nand2_1
X_0873_ _0902_/A _0879_/B vssd1 vssd1 vccd1 vccd1 _0911_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_27_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1425_ _1425_/A _1425_/B vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__nand2_1
X_1287_ _1287_/A _1287_/B vssd1 vssd1 vccd1 vccd1 _1289_/A sky130_fd_sc_hd__nand2_1
X_1356_ _1356_/A _1416_/B _1588_/B vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__and3_1
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1210_ _1210_/A _1210_/B _1237_/A vssd1 vssd1 vccd1 vccd1 _1211_/B sky130_fd_sc_hd__nand3_1
X_1072_ _0978_/B _0979_/A _0976_/Y vssd1 vssd1 vccd1 vccd1 _1073_/B sky130_fd_sc_hd__a21o_1
X_1141_ _1303_/A _1303_/B _1141_/C _1141_/D vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__or4_1
X_1635__18 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1705_/CLK sky130_fd_sc_hd__inv_2
X_0856_ _0907_/A _0856_/B vssd1 vssd1 vccd1 vccd1 _0863_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0925_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0926_/C sky130_fd_sc_hd__inv_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1408_ _1588_/B input3/X vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__and2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ _1339_/A _1339_/B _1588_/B vssd1 vssd1 vccd1 vccd1 _1340_/A sky130_fd_sc_hd__and3_1
XFILLER_0_32_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1690_ _1690_/CLK hold29/X vssd1 vssd1 vccd1 vccd1 _1690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1055_ _1055_/A vssd1 vssd1 vccd1 vccd1 _1057_/A sky130_fd_sc_hd__inv_2
X_1124_ _1124_/A _1124_/B vssd1 vssd1 vccd1 vccd1 _1178_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0839_ _1668_/Q _1678_/Q vssd1 vssd1 vccd1 vccd1 _0841_/B sky130_fd_sc_hd__nand2_1
X_0908_ _0908_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0911_/A sky130_fd_sc_hd__nand2_1
Xoutput29 _1689_/Q vssd1 vssd1 vccd1 vccd1 p[4] sky130_fd_sc_hd__buf_12
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1673_ _1673_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _1673_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1107_ _1107_/A _1667_/Q _1681_/Q vssd1 vssd1 vccd1 vccd1 _1109_/B sky130_fd_sc_hd__and3_1
X_1038_ _1669_/Q _1680_/Q vssd1 vssd1 vccd1 vccd1 _1051_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1604__43 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1675_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1725_ _1725_/CLK _1725_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
X_1587_ _1587_/A hold74/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__nand2_1
Xhold103 hold77/A vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1441_ _1441_/A _1735_/Q vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__nand2_1
X_1510_ hold36/X hold8/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__nand2_2
X_1595__34 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1666_/CLK sky130_fd_sc_hd__inv_2
X_1372_ _1376_/B _1376_/A vssd1 vssd1 vccd1 vccd1 _1374_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1708_ _1708_/CLK _1708_/D vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0941_ _1263_/C _0962_/B _0939_/C vssd1 vssd1 vccd1 vccd1 _0942_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0872_ _0872_/A _0872_/B vssd1 vssd1 vccd1 vccd1 _0879_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1355_ _1230_/A _1230_/C _1230_/B vssd1 vssd1 vccd1 vccd1 _1356_/A sky130_fd_sc_hd__a21o_1
X_1424_ hold27/X vssd1 vssd1 vccd1 vccd1 _1425_/B sky130_fd_sc_hd__inv_2
X_1286_ _1288_/B vssd1 vssd1 vccd1 vccd1 _1287_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1071_ _1071_/A _1074_/A vssd1 vssd1 vccd1 vccd1 _1073_/A sky130_fd_sc_hd__nor2b_1
X_1140_ _1668_/Q vssd1 vssd1 vccd1 vccd1 _1303_/B sky130_fd_sc_hd__inv_2
X_0924_ _1680_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _0929_/A sky130_fd_sc_hd__nand2_1
X_0855_ _0867_/B vssd1 vssd1 vccd1 vccd1 _0856_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1407_ _1407_/A vssd1 vssd1 vccd1 vccd1 _1705_/D sky130_fd_sc_hd__clkbuf_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _1338_/A _1338_/B vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__nand2_1
X_1269_ _1269_/A vssd1 vssd1 vccd1 vccd1 _1273_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1625__63 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1695_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1054_ _1131_/A _1054_/B vssd1 vssd1 vccd1 vccd1 _1059_/A sky130_fd_sc_hd__nand2_1
X_1123_ _1124_/A _1124_/B vssd1 vssd1 vccd1 vccd1 _1179_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0907_ _0907_/A _0907_/B vssd1 vssd1 vccd1 vccd1 _0930_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0838_ _1670_/Q _1676_/Q vssd1 vssd1 vccd1 vccd1 _0841_/A sky130_fd_sc_hd__nand2_1
Xoutput19 _1685_/Q vssd1 vssd1 vccd1 vccd1 p[0] sky130_fd_sc_hd__buf_12
XFILLER_0_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1672_ _1672_/CLK _1672_/D vssd1 vssd1 vccd1 vccd1 _1672_/Q sky130_fd_sc_hd__dfxtp_2
X_1106_ _1106_/A _1669_/Q _1679_/Q vssd1 vssd1 vccd1 vccd1 _1109_/A sky130_fd_sc_hd__and3_1
X_1037_ _1037_/A _1098_/A vssd1 vssd1 vccd1 vccd1 _1070_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold104 _1734_/Q vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1724_ _1724_/CLK _1724_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1586_ hold74/X _1587_/A vssd1 vssd1 vccd1 vccd1 _1588_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1652__2 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1722_/CLK sky130_fd_sc_hd__inv_2
X_1440_ _1735_/Q _1441_/A vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__or2_1
XFILLER_0_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1371_ _1369_/Y _1370_/Y _1592_/A vssd1 vssd1 vccd1 vccd1 _1722_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1707_ _1707_/CLK _1707_/D vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ hold69/X vssd1 vssd1 vccd1 vccd1 _1671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0940_ _0940_/A vssd1 vssd1 vccd1 vccd1 _1033_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0871_ _0906_/B _0871_/B vssd1 vssd1 vccd1 vccd1 _0872_/B sky130_fd_sc_hd__nand2_1
X_1423_ hold33/X _1485_/A vssd1 vssd1 vccd1 vccd1 _1425_/A sky130_fd_sc_hd__nor2_1
X_1354_ _1352_/X _1353_/Y _1592_/A vssd1 vssd1 vccd1 vccd1 _1727_/D sky130_fd_sc_hd__a21oi_1
X_1285_ _1285_/A _1326_/B vssd1 vssd1 vccd1 vccd1 _1288_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1070_ _1070_/A _1070_/B vssd1 vssd1 vccd1 vccd1 _1074_/A sky130_fd_sc_hd__nand2_1
X_0854_ _0864_/A _0865_/A vssd1 vssd1 vccd1 vccd1 _0867_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0923_ _1339_/B _0923_/B _1337_/B vssd1 vssd1 vccd1 vccd1 _0926_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1268_ _1268_/A _1268_/B vssd1 vssd1 vccd1 vccd1 _1269_/A sky130_fd_sc_hd__nand2_1
X_1406_ _1588_/B input4/X vssd1 vssd1 vccd1 vccd1 _1407_/A sky130_fd_sc_hd__and2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ _1337_/A _1337_/B vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__nand2_1
X_1199_ _1199_/A _1200_/B _1200_/A vssd1 vssd1 vccd1 vccd1 _1201_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1640__23 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1710_/CLK sky130_fd_sc_hd__inv_2
X_1122_ _1122_/A _1151_/B vssd1 vssd1 vccd1 vccd1 _1124_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ _1053_/A _1053_/B vssd1 vssd1 vccd1 vccd1 _1131_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0906_ _0906_/A _0906_/B vssd1 vssd1 vccd1 vccd1 _0908_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0837_ _0837_/A vssd1 vssd1 vccd1 vccd1 _1734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1671_ _1671_/CLK _1671_/D vssd1 vssd1 vccd1 vccd1 _1671_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1105_ _1116_/A _1116_/C vssd1 vssd1 vccd1 vccd1 _1115_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ _1036_/A _1098_/C _1036_/C vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold105 _1493_/Y vssd1 vssd1 vccd1 vccd1 _1494_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1723_ _1723_/CLK _1723_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
X_1585_ _1590_/B _1585_/B vssd1 vssd1 vccd1 vccd1 _1587_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1019_ _1019_/A _1019_/B vssd1 vssd1 vccd1 vccd1 _1094_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1370_ _1369_/B _1370_/B _1370_/C vssd1 vssd1 vccd1 vccd1 _1370_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1706_ _1706_/CLK _1706_/D vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1568_/A _1588_/B hold68/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__and3_1
X_1499_ _1499_/A hold70/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0870_ _0870_/A _0870_/B vssd1 vssd1 vccd1 vccd1 _0906_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1422_ hold30/X _1422_/B vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__or2_1
X_1353_ _1353_/A _1353_/B vssd1 vssd1 vccd1 vccd1 _1353_/Y sky130_fd_sc_hd__nand2_1
X_1284_ _1284_/A _1310_/A _1284_/C vssd1 vssd1 vccd1 vccd1 _1326_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0999_ _0999_/A _0999_/B vssd1 vssd1 vccd1 vccd1 _1000_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0853_ _0864_/A _0865_/A vssd1 vssd1 vccd1 vccd1 _0907_/A sky130_fd_sc_hd__nor2_1
X_0922_ _0922_/A _0930_/A _0922_/C vssd1 vssd1 vccd1 vccd1 _0985_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1405_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1198_ _1240_/B _1240_/A vssd1 vssd1 vccd1 vccd1 _1200_/B sky130_fd_sc_hd__xnor2_1
X_1267_ _1273_/A vssd1 vssd1 vccd1 vccd1 _1267_/Y sky130_fd_sc_hd__inv_2
Xinput1 a[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_1336_ _1336_/A vssd1 vssd1 vccd1 vccd1 _1732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1052_ _1052_/A vssd1 vssd1 vccd1 vccd1 _1053_/B sky130_fd_sc_hd__inv_2
X_1121_ _1136_/A _1121_/B _1121_/C vssd1 vssd1 vccd1 vccd1 _1151_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1616__54 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1686_/CLK sky130_fd_sc_hd__inv_2
X_0836_ _1588_/B _1682_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _0837_/A sky130_fd_sc_hd__and3_1
X_0905_ _0905_/A _0905_/B vssd1 vssd1 vccd1 vccd1 _0926_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1319_ _1320_/B _1320_/A vssd1 vssd1 vccd1 vccd1 _1321_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1670_ _1670_/CLK _1670_/D vssd1 vssd1 vccd1 vccd1 _1670_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1104_ _1104_/A _1171_/A vssd1 vssd1 vccd1 vccd1 _1124_/A sky130_fd_sc_hd__nand2_1
X_1035_ _1036_/A _1098_/C _1036_/C vssd1 vssd1 vccd1 vccd1 _1037_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1610__49 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1681_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1584_ _1584_/A vssd1 vssd1 vccd1 vccd1 _1590_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold106 _1494_/X vssd1 vssd1 vccd1 vccd1 _1495_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1722_ _1722_/CLK _1722_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1018_ _1154_/B _1018_/B vssd1 vssd1 vccd1 vccd1 _1019_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1705_ _1705_/CLK _1705_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1567_ _1567_/A hold67/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__nand2_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ hold70/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1500_/A sky130_fd_sc_hd__or2_1
XFILLER_0_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1421_ _1492_/B _1421_/B vssd1 vssd1 vccd1 vccd1 _1422_/B sky130_fd_sc_hd__nand2_1
X_1352_ _1353_/B _1353_/A vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__or2_1
X_1283_ _1284_/A _1310_/A _1284_/C vssd1 vssd1 vccd1 vccd1 _1285_/A sky130_fd_sc_hd__a21o_1
X_1661__11 _1613_/A vssd1 vssd1 vccd1 vccd1 _1731_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_25_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0998_ _0998_/A vssd1 vssd1 vccd1 vccd1 _1341_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0922_/C sky130_fd_sc_hd__inv_2
X_0852_ _1680_/Q _1673_/Q vssd1 vssd1 vccd1 vccd1 _0865_/A sky130_fd_sc_hd__nand2_1
X_1404_ _1588_/B input5/X vssd1 vssd1 vccd1 vccd1 _1405_/A sky130_fd_sc_hd__and2_1
X_1335_ _1338_/B _1588_/B _1335_/C vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__and3_1
X_1197_ _1197_/A _1197_/B vssd1 vssd1 vccd1 vccd1 _1240_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1266_ _1268_/A _1268_/B vssd1 vssd1 vccd1 vccd1 _1273_/A sky130_fd_sc_hd__nor2_1
Xinput2 a[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1051_ _1051_/A vssd1 vssd1 vccd1 vccd1 _1053_/A sky130_fd_sc_hd__inv_2
X_1120_ _1196_/A vssd1 vssd1 vccd1 vccd1 _1121_/C sky130_fd_sc_hd__inv_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0904_ _0923_/B vssd1 vssd1 vccd1 vccd1 _0905_/B sky130_fd_sc_hd__inv_2
X_0835_ _0835_/A vssd1 vssd1 vccd1 vccd1 _1735_/D sky130_fd_sc_hd__clkbuf_1
X_1631__69 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ _1318_/A _1318_/B vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__nand2_1
X_1249_ _1249_/A _1249_/B vssd1 vssd1 vccd1 vccd1 _1250_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1103_ _1158_/A _1103_/B _1103_/C vssd1 vssd1 vccd1 vccd1 _1171_/A sky130_fd_sc_hd__nand3_2
X_1034_ _1034_/A _1094_/C _1034_/C vssd1 vssd1 vccd1 vccd1 _1098_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1721_ _1721_/CLK _1721_/D vssd1 vssd1 vccd1 vccd1 _1721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1583_ hold38/X _1583_/B vssd1 vssd1 vccd1 vccd1 _1584_/A sky130_fd_sc_hd__and2b_1
Xhold107 _1721_/Q vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1017_ _1027_/B vssd1 vssd1 vccd1 vccd1 _1018_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1704_ _1704_/CLK _1704_/D vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1566_ hold67/X _1567_/A vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__or2_1
X_1497_ _1506_/A _1497_/B vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__nor2_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1420_ hold99/X vssd1 vssd1 vccd1 vccd1 _1421_/B sky130_fd_sc_hd__inv_2
X_1351_ _1351_/A _1351_/B vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__nand2_1
X_1282_ _1317_/A vssd1 vssd1 vccd1 vccd1 _1284_/C sky130_fd_sc_hd__inv_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ _0997_/A _0997_/B vssd1 vssd1 vccd1 vccd1 _0998_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1549_ hold92/X _1549_/B vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__nor2_1
X_1637__20 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ _0920_/A _0921_/A vssd1 vssd1 vccd1 vccd1 _0985_/A sky130_fd_sc_hd__nand2_1
X_0851_ _1679_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _0864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1265_ _1307_/B _1265_/B vssd1 vssd1 vccd1 vccd1 _1268_/B sky130_fd_sc_hd__nand2_1
X_1403_ _1403_/A vssd1 vssd1 vccd1 vccd1 _1707_/D sky130_fd_sc_hd__clkbuf_1
X_1334_ _1334_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1335_/C sky130_fd_sc_hd__nand2_1
X_1196_ _1196_/A _1667_/Q _1679_/Q vssd1 vssd1 vccd1 vccd1 _1240_/B sky130_fd_sc_hd__and3_1
Xinput3 a[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1050_ _1050_/A _1050_/B vssd1 vssd1 vccd1 vccd1 _1112_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0834_ _1588_/B _0834_/B vssd1 vssd1 vccd1 vccd1 _0835_/A sky130_fd_sc_hd__and2_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0903_ _0903_/A _0909_/A vssd1 vssd1 vccd1 vccd1 _0923_/B sky130_fd_sc_hd__nand2_1
X_1248_ _1248_/A _1248_/B vssd1 vssd1 vccd1 vccd1 _1249_/B sky130_fd_sc_hd__xnor2_1
X_1317_ _1317_/A _1667_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1320_/B sky130_fd_sc_hd__and3_1
X_1179_ _1179_/A vssd1 vssd1 vccd1 vccd1 _1180_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1655__5 _1613_/A vssd1 vssd1 vccd1 vccd1 _1725_/CLK sky130_fd_sc_hd__inv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__0832_ clkbuf_0__0832_/X vssd1 vssd1 vccd1 vccd1 _1630__68/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ _1187_/A vssd1 vssd1 vccd1 vccd1 _1103_/C sky130_fd_sc_hd__inv_2
X_1033_ _1033_/A _1033_/B vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1720_ _1720_/CLK _1720_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1582_ hold73/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1024_/A _1025_/A vssd1 vssd1 vccd1 vccd1 _1027_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1703_ _1703_/CLK _1703_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1570_/A _1585_/B vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__nand2_1
X_1496_ hold5/X _1496_/B vssd1 vssd1 vccd1 vccd1 _1497_/B sky130_fd_sc_hd__nor2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1350_ _1350_/A vssd1 vssd1 vccd1 vccd1 _1728_/D sky130_fd_sc_hd__inv_2
X_1281_ _1668_/Q _1676_/Q vssd1 vssd1 vccd1 vccd1 _1317_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0996_ _0926_/A _0926_/B _0926_/C vssd1 vssd1 vccd1 vccd1 _0997_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_41_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1479_ _1479_/A hold80/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__nand2_1
X_1548_ hold36/A vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0850_ _1293_/A _0850_/B vssd1 vssd1 vccd1 vccd1 _1218_/B sky130_fd_sc_hd__nand2_1
X_1402_ _1588_/B input6/X vssd1 vssd1 vccd1 vccd1 _1403_/A sky130_fd_sc_hd__and2_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1264_ _1667_/Q _1678_/Q _1668_/Q _1677_/Q vssd1 vssd1 vccd1 vccd1 _1265_/B sky130_fd_sc_hd__a22o_1
Xinput4 a[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_1333_ _1333_/A vssd1 vssd1 vccd1 vccd1 _1338_/B sky130_fd_sc_hd__inv_2
X_1195_ _1246_/A vssd1 vssd1 vccd1 vccd1 _1203_/A sky130_fd_sc_hd__inv_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0979_ _0979_/A _0979_/B vssd1 vssd1 vccd1 vccd1 _0981_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0902_ _0902_/A _0911_/B vssd1 vssd1 vccd1 vccd1 _0909_/A sky130_fd_sc_hd__or2_1
X_0833_ _1700_/Q vssd1 vssd1 vccd1 vccd1 _1588_/B sky130_fd_sc_hd__inv_8
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1247_ _1210_/A _1237_/A _1246_/Y vssd1 vssd1 vccd1 vccd1 _1249_/A sky130_fd_sc_hd__a21oi_1
X_1178_ _1178_/A _1178_/B vssd1 vssd1 vccd1 vccd1 _1180_/A sky130_fd_sc_hd__nand2_1
X_1316_ _1326_/B _1326_/A vssd1 vssd1 vccd1 vccd1 _1327_/A sky130_fd_sc_hd__or2_1
X_1607__46 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1678_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0831_ clkbuf_0__0831_/X vssd1 vssd1 vccd1 vccd1 _1612__51/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1101_ _1101_/A _1187_/A vssd1 vssd1 vccd1 vccd1 _1104_/A sky130_fd_sc_hd__nand2_1
X_1032_ _1034_/A _1094_/C vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1581_ hold40/X vssd1 vssd1 vccd1 vccd1 _1669_/D sky130_fd_sc_hd__clkbuf_1
X_1598__37 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1669_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1015_ _1024_/A _1025_/A vssd1 vssd1 vccd1 vccd1 _1154_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ _1702_/CLK _1702_/D vssd1 vssd1 vccd1 vccd1 _1702_/Q sky130_fd_sc_hd__dfxtp_1
X_1564_ _1577_/A vssd1 vssd1 vccd1 vccd1 _1585_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1495_/A vssd1 vssd1 vccd1 vccd1 _1687_/D sky130_fd_sc_hd__clkbuf_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1280_ _1280_/A _1280_/B vssd1 vssd1 vccd1 vccd1 _1310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0995_ _0995_/A _0995_/B _0995_/C vssd1 vssd1 vccd1 vccd1 _1004_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1547_ _1547_/A vssd1 vssd1 vccd1 vccd1 _1676_/D sky130_fd_sc_hd__clkbuf_1
X_1478_ hold80/X _1479_/A vssd1 vssd1 vccd1 vccd1 _1480_/A sky130_fd_sc_hd__or2_1
X_1628__66 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1698_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1401_ _1401_/A vssd1 vssd1 vccd1 vccd1 _1708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1194_ _1194_/A _1239_/A vssd1 vssd1 vccd1 vccd1 _1246_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1263_ _1303_/A _1303_/B _1263_/C _1263_/D vssd1 vssd1 vccd1 vccd1 _1307_/B sky130_fd_sc_hd__or4_1
Xinput5 a[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_1332_ _1329_/Y _1330_/X _1592_/A vssd1 vssd1 vccd1 vccd1 _1733_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ _0976_/Y _0978_/B vssd1 vssd1 vccd1 vccd1 _0979_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0901_ _0901_/A _0911_/B _0902_/A vssd1 vssd1 vccd1 vccd1 _0903_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1315_ _1315_/A _1323_/A vssd1 vssd1 vccd1 vccd1 _1326_/A sky130_fd_sc_hd__nand2_1
X_1246_ _1246_/A _1246_/B vssd1 vssd1 vccd1 vccd1 _1246_/Y sky130_fd_sc_hd__nor2_1
X_1177_ _1209_/B _1208_/A vssd1 vssd1 vccd1 vccd1 _1182_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0830_ clkbuf_0__0830_/X vssd1 vssd1 vccd1 vccd1 _1659__9/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1031_ _1094_/B _1031_/B _1031_/C vssd1 vssd1 vccd1 vccd1 _1094_/C sky130_fd_sc_hd__nand3_2
X_1100_ _1672_/Q _1676_/Q vssd1 vssd1 vccd1 vccd1 _1187_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1229_ _1229_/A _1229_/B _1229_/C vssd1 vssd1 vccd1 vccd1 _1230_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1580_ _1580_/A _1588_/B hold39/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__and3_1
XFILLER_0_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ _1671_/Q _1678_/Q vssd1 vssd1 vccd1 vccd1 _1025_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_0__0832_ _1613_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0832_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1701_ _1701_/CLK _1701_/D vssd1 vssd1 vccd1 vccd1 _1701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1563_ _1563_/A hold95/A vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__nand2_1
X_1632_ _1632_/A vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__buf_1
X_1494_ _1494_/A _1588_/B _1494_/C vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__and3_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0994_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0995_/C sky130_fd_sc_hd__inv_2
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1477_ hold89/X vssd1 vssd1 vccd1 vccd1 _1479_/A sky130_fd_sc_hd__inv_2
X_1546_ _1546_/A _1588_/B _1546_/C vssd1 vssd1 vccd1 vccd1 _1547_/A sky130_fd_sc_hd__and3_1
X_1643__26 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1400_ _1588_/B input7/X vssd1 vssd1 vccd1 vccd1 _1401_/A sky130_fd_sc_hd__and2_1
X_1331_ _1700_/Q vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1193_ _1193_/A _1193_/B vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__or2_1
XFILLER_0_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1262_ _1307_/A _1262_/B vssd1 vssd1 vccd1 vccd1 _1268_/A sky130_fd_sc_hd__nand2_1
Xinput6 a[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ _0977_/A _0977_/B vssd1 vssd1 vccd1 vccd1 _0978_/B sky130_fd_sc_hd__nand2_1
X_1529_ _1529_/A hold60/A vssd1 vssd1 vccd1 vccd1 _1534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0900_ _0909_/B _0900_/B vssd1 vssd1 vccd1 vccd1 _0911_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1314_ _1314_/A _1314_/B vssd1 vssd1 vccd1 vccd1 _1323_/A sky130_fd_sc_hd__nand2_1
X_1245_ _1245_/A _1245_/B vssd1 vssd1 vccd1 vccd1 _1250_/A sky130_fd_sc_hd__nand2_1
X_1176_ _1176_/A _1176_/B vssd1 vssd1 vccd1 vccd1 _1208_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1030_ _1159_/A _1030_/B vssd1 vssd1 vccd1 vccd1 _1034_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1612__51 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1683_/CLK sky130_fd_sc_hd__inv_2
X_1228_ _1228_/A _1232_/A vssd1 vssd1 vccd1 vccd1 _1414_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1159_ _1159_/A _1159_/B _1159_/C vssd1 vssd1 vccd1 vccd1 _1188_/A sky130_fd_sc_hd__or3_2
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _1677_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _1024_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_0__0831_ _1594_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0831_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1700_ _1632_/A _1700_/D vssd1 vssd1 vccd1 vccd1 _1700_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ hold66/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__inv_2
X_1493_ _1492_/B _1506_/A _1492_/A vssd1 vssd1 vccd1 vccd1 _1493_/Y sky130_fd_sc_hd__o21ai_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1649__32 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1719_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0993_ _0993_/A _0994_/A vssd1 vssd1 vccd1 vccd1 _1003_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1476_ _1476_/A hold88/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__nand2_1
X_1545_ _1545_/A hold93/X vssd1 vssd1 vccd1 vccd1 _1546_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1658__8 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1728_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1261_ _1669_/Q _1676_/Q _1670_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1262_/B sky130_fd_sc_hd__a22o_1
X_1330_ _1330_/A _1330_/B _1330_/C vssd1 vssd1 vccd1 vccd1 _1330_/X sky130_fd_sc_hd__and3_1
X_1192_ _1192_/A _1193_/B _1193_/A vssd1 vssd1 vccd1 vccd1 _1194_/A sky130_fd_sc_hd__nand3_1
X_1619__57 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1689_/CLK sky130_fd_sc_hd__inv_2
Xinput7 a[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ _0977_/B _0977_/A vssd1 vssd1 vccd1 vccd1 _0976_/Y sky130_fd_sc_hd__nor2_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1459_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1461_/A sky130_fd_sc_hd__inv_2
X_1528_ _1528_/A vssd1 vssd1 vccd1 vccd1 _1529_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1244_ _1244_/A _1244_/B vssd1 vssd1 vccd1 vccd1 _1245_/B sky130_fd_sc_hd__nand2_1
X_1313_ _1314_/B _1314_/A vssd1 vssd1 vccd1 vccd1 _1315_/A sky130_fd_sc_hd__or2_1
X_1175_ _1175_/A vssd1 vssd1 vccd1 vccd1 _1209_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0959_ _1031_/C vssd1 vssd1 vccd1 vccd1 _1030_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 b[1] vssd1 vssd1 vccd1 vccd1 _1394_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1158_ _1158_/A _1158_/B vssd1 vssd1 vccd1 vccd1 _1168_/A sky130_fd_sc_hd__nand2_1
X_1227_ _1276_/B _1227_/B vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__nand2_1
X_1089_ _1089_/A _1671_/Q _1677_/Q vssd1 vssd1 vccd1 vccd1 _1091_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1012_ _1154_/A _1012_/B vssd1 vssd1 vccd1 vccd1 _1019_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__0830_ _1593_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0830_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1492_/A _1492_/B _1506_/A vssd1 vssd1 vccd1 vccd1 _1494_/A sky130_fd_sc_hd__or3_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1561_/A vssd1 vssd1 vccd1 vccd1 _1672_/D sky130_fd_sc_hd__clkbuf_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664__14 _1613_/A vssd1 vssd1 vccd1 vccd1 _1734_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0992_ _0992_/A _0992_/B vssd1 vssd1 vccd1 vccd1 _0994_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1613_ _1613_/A vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__buf_1
XFILLER_0_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1544_ hold93/X _1545_/A vssd1 vssd1 vccd1 vccd1 _1546_/A sky130_fd_sc_hd__or2_1
X_1475_ hold50/X _1474_/X _1588_/B vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__o21a_1
XFILLER_0_32_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1191_ _1191_/A _1239_/C vssd1 vssd1 vccd1 vccd1 _1193_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1260_ _1260_/A _1260_/B _1303_/C _1303_/D vssd1 vssd1 vccd1 vccd1 _1307_/A sky130_fd_sc_hd__or4_1
Xinput8 a[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1634__17 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1704_/CLK sky130_fd_sc_hd__inv_2
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ _1067_/C _0975_/B vssd1 vssd1 vccd1 vccd1 _0977_/A sky130_fd_sc_hd__nand2b_1
X_1527_ hold62/X vssd1 vssd1 vccd1 vccd1 _1679_/D sky130_fd_sc_hd__clkbuf_1
X_1389_ _1389_/A vssd1 vssd1 vccd1 vccd1 _1714_/D sky130_fd_sc_hd__clkbuf_1
X_1458_ _1458_/A hold88/A vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__nand2_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1174_ _1176_/B _1176_/A vssd1 vssd1 vccd1 vccd1 _1175_/A sky130_fd_sc_hd__nor2_1
X_1243_ _1248_/B _1248_/A vssd1 vssd1 vccd1 vccd1 _1244_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1312_ _1312_/A vssd1 vssd1 vccd1 vccd1 _1314_/A sky130_fd_sc_hd__inv_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0958_ _1088_/A _1089_/A vssd1 vssd1 vccd1 vccd1 _1031_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0889_ _1681_/Q vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__inv_2
XFILLER_0_27_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 b[2] vssd1 vssd1 vccd1 vccd1 _1392_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1632_/A sky130_fd_sc_hd__clkbuf_16
X_1157_ _1157_/A vssd1 vssd1 vccd1 vccd1 _1158_/B sky130_fd_sc_hd__inv_2
X_1226_ _1669_/Q _1678_/Q _1670_/Q _1677_/Q vssd1 vssd1 vccd1 vccd1 _1227_/B sky130_fd_sc_hd__a22o_1
X_1088_ _1088_/A _1673_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1091_/A sky130_fd_sc_hd__and3_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1603__42 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1674_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _1023_/B vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ _1209_/A _1209_/B vssd1 vssd1 vccd1 vccd1 _1210_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1560_ _1560_/A _1588_/B _1560_/C vssd1 vssd1 vccd1 vccd1 _1561_/A sky130_fd_sc_hd__and3_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1489_/X hold31/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__a21oi_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1689_ _1689_/CLK hold35/X vssd1 vssd1 vccd1 vccd1 _1689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0991_ _0991_/A _1000_/A vssd1 vssd1 vccd1 vccd1 _0992_/B sky130_fd_sc_hd__nand2_1
X_1474_ hold49/X hold81/A _1471_/A vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__o21ba_1
X_1543_ _1549_/B _1543_/B vssd1 vssd1 vccd1 vccd1 _1545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1190_ _1190_/A _1190_/B vssd1 vssd1 vccd1 vccd1 _1239_/C sky130_fd_sc_hd__nand2_1
Xinput9 b[0] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0974_ _0974_/A _0974_/B vssd1 vssd1 vccd1 vccd1 _0975_/B sky130_fd_sc_hd__nand2_1
X_1457_ hold57/X _1456_/X _1588_/B vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__o21a_1
X_1526_ _1526_/A _1588_/B hold61/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__and3_1
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1388_ _1588_/B _1388_/B vssd1 vssd1 vccd1 vccd1 _1389_/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1624__62 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1694_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1311_ _1318_/A _1311_/B vssd1 vssd1 vccd1 vccd1 _1312_/A sky130_fd_sc_hd__nand2_1
X_1242_ _1248_/A _1248_/B vssd1 vssd1 vccd1 vccd1 _1244_/A sky130_fd_sc_hd__nand2b_1
X_1173_ _1173_/A _1192_/A vssd1 vssd1 vccd1 vccd1 _1176_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0957_ _1678_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _1089_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0888_ _0888_/A _0888_/B vssd1 vssd1 vccd1 vccd1 _1334_/B sky130_fd_sc_hd__nand2_1
X_1509_ _1592_/A _1511_/B vssd1 vssd1 vccd1 vccd1 _1682_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_18_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 b[3] vssd1 vssd1 vccd1 vccd1 _1390_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1156_ _1156_/A _1156_/B _1159_/B vssd1 vssd1 vccd1 vccd1 _1157_/A sky130_fd_sc_hd__nand3_1
X_1087_ _1098_/A _1098_/C vssd1 vssd1 vccd1 vccd1 _1097_/A sky130_fd_sc_hd__nand2_1
X_1225_ _1260_/A _1260_/B _1263_/C _1263_/D vssd1 vssd1 vccd1 vccd1 _1276_/B sky130_fd_sc_hd__or4_1
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ _1020_/A _1021_/A vssd1 vssd1 vccd1 vccd1 _1023_/B sky130_fd_sc_hd__nand2_1
X_1208_ _1208_/A _1208_/B vssd1 vssd1 vccd1 vccd1 _1209_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ _1667_/Q vssd1 vssd1 vccd1 vccd1 _1303_/A sky130_fd_sc_hd__inv_2
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1490_ _1506_/A hold30/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__nand2_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1688_ _1688_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 _1688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0990_ _1000_/A _0991_/A vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1473_ hold49/X hold88/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__nor2_1
X_1542_ _1542_/A vssd1 vssd1 vccd1 vccd1 _1549_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ _0974_/B _0974_/A vssd1 vssd1 vccd1 vccd1 _1067_/C sky130_fd_sc_hd__nor2_1
X_1387_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1715_/D sky130_fd_sc_hd__clkbuf_1
X_1456_ hold56/X _1434_/A _1453_/A vssd1 vssd1 vccd1 vccd1 _1456_/X sky130_fd_sc_hd__o21ba_1
X_1525_ _1525_/A hold60/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1241_ _1241_/A _1241_/B _1241_/C vssd1 vssd1 vccd1 vccd1 _1248_/B sky130_fd_sc_hd__and3_1
X_1310_ _1310_/A _1310_/B vssd1 vssd1 vccd1 vccd1 _1311_/B sky130_fd_sc_hd__nand2_1
X_1172_ _1172_/A _1193_/A _1172_/C vssd1 vssd1 vccd1 vccd1 _1192_/A sky130_fd_sc_hd__nand3_1
X_0956_ _1676_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _1088_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0887_ _0895_/A _0896_/A vssd1 vssd1 vccd1 vccd1 _0888_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1439_ hold86/X vssd1 vssd1 vccd1 vccd1 _1441_/A sky130_fd_sc_hd__inv_2
X_1508_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1511_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 b[4] vssd1 vssd1 vccd1 vccd1 _1388_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1224_ _1670_/Q vssd1 vssd1 vccd1 vccd1 _1260_/B sky130_fd_sc_hd__inv_2
X_1155_ _1155_/A _1188_/B vssd1 vssd1 vccd1 vccd1 _1159_/B sky130_fd_sc_hd__nand2_1
X_1086_ _1074_/A _1073_/B _1071_/A vssd1 vssd1 vccd1 vccd1 _1178_/A sky130_fd_sc_hd__a21o_1
X_0939_ _1263_/C _0962_/B _0939_/C vssd1 vssd1 vccd1 vccd1 _0940_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ _1207_/A _1207_/B vssd1 vssd1 vccd1 vccd1 _1211_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ _1150_/A _1197_/A vssd1 vssd1 vccd1 vccd1 _1149_/A sky130_fd_sc_hd__nand2_1
X_1069_ _1070_/A _1070_/B vssd1 vssd1 vccd1 vccd1 _1071_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1687_ _1687_/CLK _1687_/D vssd1 vssd1 vccd1 vccd1 _1687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1472_ _1470_/X hold19/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__a21oi_1
X_1541_ hold41/X _1541_/B vssd1 vssd1 vccd1 vccd1 _1542_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ _0972_/A _1260_/A _0999_/B vssd1 vssd1 vccd1 vccd1 _0974_/A sky130_fd_sc_hd__or3b_1
X_1524_ hold60/X _1525_/A vssd1 vssd1 vccd1 vccd1 _1526_/A sky130_fd_sc_hd__or2_1
X_1386_ _1588_/B _1386_/B vssd1 vssd1 vccd1 vccd1 _1387_/A sky130_fd_sc_hd__and2_1
X_1455_ hold56/X hold88/A vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1240_ _1240_/A _1240_/B vssd1 vssd1 vccd1 vccd1 _1241_/C sky130_fd_sc_hd__nand2_1
X_1171_ _1171_/A vssd1 vssd1 vccd1 vccd1 _1172_/C sky130_fd_sc_hd__inv_2
X_0955_ _0955_/A vssd1 vssd1 vccd1 vccd1 _0979_/A sky130_fd_sc_hd__inv_2
X_1615__53 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1685_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ _0886_/A _0901_/A _0891_/C vssd1 vssd1 vccd1 vccd1 _1337_/B sky130_fd_sc_hd__nand3_2
X_1507_ hold84/X _1506_/Y _1592_/A vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1438_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1496_/B sky130_fd_sc_hd__inv_2
X_1369_ _1369_/A _1369_/B vssd1 vssd1 vccd1 vccd1 _1369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 b[5] vssd1 vssd1 vccd1 vccd1 _1386_/B sky130_fd_sc_hd__clkbuf_1
X_1154_ _1154_/A _1154_/B vssd1 vssd1 vccd1 vccd1 _1188_/B sky130_fd_sc_hd__nand2_1
X_1223_ _1233_/A _1233_/B vssd1 vssd1 vccd1 vccd1 _1228_/A sky130_fd_sc_hd__nand2_1
X_1085_ _1229_/A _1229_/C vssd1 vssd1 vccd1 vccd1 _1252_/B sky130_fd_sc_hd__nand2_2
X_0938_ _1677_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _0939_/C sky130_fd_sc_hd__nand2_1
X_0869_ _0869_/A vssd1 vssd1 vccd1 vccd1 _0870_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1137_ _1137_/A _1137_/B _1137_/C vssd1 vssd1 vccd1 vccd1 _1197_/A sky130_fd_sc_hd__or3_2
X_1206_ _1208_/A _1208_/B _1175_/A vssd1 vssd1 vccd1 vccd1 _1207_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1068_ _1068_/A _1116_/A vssd1 vssd1 vccd1 vccd1 _1070_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1686_ _1686_/CLK _1686_/D vssd1 vssd1 vccd1 vccd1 _1686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1646__29 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1716_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1540_ hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__inv_2
X_1471_ _1471_/A hold18/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__nand2_1
X_1660__10 _1613_/A vssd1 vssd1 vccd1 vccd1 _1730_/CLK sky130_fd_sc_hd__inv_2
X_1669_ _1669_/CLK _1669_/D vssd1 vssd1 vccd1 vccd1 _1669_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0832_ clkbuf_0__0832_/X vssd1 vssd1 vccd1 vccd1 _1631__69/A sky130_fd_sc_hd__clkbuf_16
X_0971_ _1061_/B _0971_/B vssd1 vssd1 vccd1 vccd1 _0974_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1454_ _1452_/X hold22/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__a21oi_1
X_1523_ _1528_/A _1543_/B vssd1 vssd1 vccd1 vccd1 _1525_/A sky130_fd_sc_hd__nand2_1
X_1385_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1170_ _1170_/A _1171_/A vssd1 vssd1 vccd1 vccd1 _1173_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0954_ _0989_/B _0988_/A _0953_/Y vssd1 vssd1 vccd1 vccd1 _0955_/A sky130_fd_sc_hd__a21oi_1
X_1630__68 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1701_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0885_ _0885_/A _1359_/A vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1506_ _1506_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _1506_/Y sky130_fd_sc_hd__nand2_1
X_1437_ hold24/X _1437_/B vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__nor2_1
X_1299_ _1299_/A vssd1 vssd1 vccd1 vccd1 _1299_/Y sky130_fd_sc_hd__inv_2
X_1368_ _1370_/B _1370_/C vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 b[6] vssd1 vssd1 vccd1 vccd1 _1384_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1153_ _1153_/A _1153_/B vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__nand2_1
X_1222_ _1230_/A _1222_/B vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__nand2_1
X_1084_ _1351_/B _1083_/Y _1080_/A vssd1 vssd1 vccd1 vccd1 _1229_/C sky130_fd_sc_hd__o21a_1
X_0937_ _1678_/Q vssd1 vssd1 vccd1 vccd1 _1263_/C sky130_fd_sc_hd__inv_2
X_0868_ _0868_/A vssd1 vssd1 vccd1 vccd1 _0870_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1136_ _1136_/A _1136_/B vssd1 vssd1 vccd1 vccd1 _1150_/A sky130_fd_sc_hd__nand2_1
X_1205_ _1210_/B _1237_/A vssd1 vssd1 vccd1 vccd1 _1207_/A sky130_fd_sc_hd__nand2_1
X_1067_ _1067_/A _1116_/C _1067_/C vssd1 vssd1 vccd1 vccd1 _1116_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1685_ _1685_/CLK _1685_/D vssd1 vssd1 vccd1 vccd1 _1685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1119_ _1119_/A _1196_/A vssd1 vssd1 vccd1 vccd1 _1122_/A sky130_fd_sc_hd__nand2_1
X_1653__3 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1723_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_34_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1470_ hold18/X _1471_/A vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1668_ _1668_/CLK _1668_/D vssd1 vssd1 vccd1 vccd1 _1668_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__0831_ clkbuf_0__0831_/X vssd1 vssd1 vccd1 vccd1 _1611__50/A sky130_fd_sc_hd__clkbuf_16
X_0970_ _1106_/A _1107_/A vssd1 vssd1 vccd1 vccd1 _0971_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1453_ _1453_/A hold21/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__nand2_1
X_1522_ hold37/A vssd1 vssd1 vccd1 vccd1 _1543_/B sky130_fd_sc_hd__inv_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1384_ _1588_/B _1384_/B vssd1 vssd1 vccd1 vccd1 _1385_/A sky130_fd_sc_hd__and2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0953_ _0953_/A _0953_/B vssd1 vssd1 vccd1 vccd1 _0953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0884_ _0891_/C vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__inv_2
X_1505_ _1431_/B hold83/X _1461_/A vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1436_ _1436_/A vssd1 vssd1 vccd1 vccd1 _1437_/B sky130_fd_sc_hd__inv_2
X_1367_ _1367_/A vssd1 vssd1 vccd1 vccd1 _1723_/D sky130_fd_sc_hd__clkbuf_1
X_1298_ _1361_/B _1301_/A vssd1 vssd1 vccd1 vccd1 _1302_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 b[7] vssd1 vssd1 vccd1 vccd1 _1382_/B sky130_fd_sc_hd__clkbuf_1
X_1221_ _1221_/A _1221_/B vssd1 vssd1 vccd1 vccd1 _1222_/B sky130_fd_sc_hd__nand2_1
X_1152_ _1199_/A _1152_/B vssd1 vssd1 vccd1 vccd1 _1176_/B sky130_fd_sc_hd__nand2_1
X_1083_ _1083_/A vssd1 vssd1 vccd1 vccd1 _1083_/Y sky130_fd_sc_hd__inv_2
X_0936_ _0982_/A _0982_/B vssd1 vssd1 vccd1 vccd1 _0980_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0867_ _0906_/A _0867_/B vssd1 vssd1 vccd1 vccd1 _0872_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1419_ hold16/X hold96/X vssd1 vssd1 vccd1 vccd1 _1492_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1600__39 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1671_/CLK sky130_fd_sc_hd__inv_2
X_1204_ _1246_/A _1246_/B vssd1 vssd1 vccd1 vccd1 _1237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1135_ _1135_/A vssd1 vssd1 vccd1 vccd1 _1136_/B sky130_fd_sc_hd__inv_2
X_1066_ _1067_/A _1116_/C _1067_/C vssd1 vssd1 vccd1 vccd1 _1068_/A sky130_fd_sc_hd__a21o_1
X_0919_ _1079_/C _0919_/B vssd1 vssd1 vccd1 vccd1 _0921_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1684_ _1684_/CLK _1684_/D vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1049_ _1132_/B _1049_/B vssd1 vssd1 vccd1 vccd1 _1050_/B sky130_fd_sc_hd__nor2_1
X_1118_ _1668_/Q _1680_/Q vssd1 vssd1 vccd1 vccd1 _1196_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1667_ _1667_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _1667_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__0830_ clkbuf_0__0830_/X vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1383_ _1383_/A vssd1 vssd1 vccd1 vccd1 _1717_/D sky130_fd_sc_hd__clkbuf_1
X_1452_ hold21/X _1453_/A vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__or2_1
X_1521_ _1521_/A hold64/A vssd1 vssd1 vccd1 vccd1 _1528_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1719_ _1719_/CLK _1719_/D vssd1 vssd1 vccd1 vccd1 _1719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ _0999_/A _0999_/B vssd1 vssd1 vccd1 vccd1 _0988_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1504_ _1504_/A vssd1 vssd1 vccd1 vccd1 _1684_/D sky130_fd_sc_hd__clkbuf_1
X_0883_ _1358_/A _1358_/B vssd1 vssd1 vccd1 vccd1 _0891_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1435_ hold21/X _1451_/A vssd1 vssd1 vccd1 vccd1 _1436_/A sky130_fd_sc_hd__nor2_1
X_1366_ _1366_/A _1370_/B _1588_/B vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__and3_1
X_1297_ _1369_/B _1364_/B vssd1 vssd1 vccd1 vccd1 _1301_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1621__59 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1691_/CLK sky130_fd_sc_hd__inv_2
X_1606__45 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1677_/CLK sky130_fd_sc_hd__inv_2
Xinput17 control vssd1 vssd1 vccd1 vccd1 _1503_/B sky130_fd_sc_hd__clkbuf_1
X_1151_ _1151_/A _1151_/B _1151_/C vssd1 vssd1 vccd1 vccd1 _1152_/B sky130_fd_sc_hd__nand3_1
X_1220_ _1252_/B _1220_/B vssd1 vssd1 vccd1 vccd1 _1230_/A sky130_fd_sc_hd__nand2_1
X_1082_ _1347_/A _1347_/B _1082_/C vssd1 vssd1 vccd1 vccd1 _1229_/A sky130_fd_sc_hd__nand3_2
X_0866_ _0866_/A _0866_/B vssd1 vssd1 vccd1 vccd1 _0906_/A sky130_fd_sc_hd__nand2_1
X_0935_ _0935_/A _0985_/B vssd1 vssd1 vccd1 vccd1 _0982_/B sky130_fd_sc_hd__or2_1
XFILLER_0_15_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1418_ _1418_/A vssd1 vssd1 vccd1 vccd1 _1701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1349_ _0984_/A _1004_/B _1345_/B _1348_/Y vssd1 vssd1 vccd1 vccd1 _1350_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1597__36 _1612__51/A vssd1 vssd1 vccd1 vccd1 _1668_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1134_ _1134_/A _1134_/B _1137_/B vssd1 vssd1 vccd1 vccd1 _1135_/A sky130_fd_sc_hd__nand3_1
X_1203_ _1203_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1210_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1065_ _1065_/A _1112_/C _1065_/C vssd1 vssd1 vccd1 vccd1 _1116_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0849_ _0849_/A _0849_/B vssd1 vssd1 vccd1 vccd1 _0850_/B sky130_fd_sc_hd__nand2_1
X_0918_ _1680_/Q _1671_/Q _1679_/Q _1672_/Q vssd1 vssd1 vccd1 vccd1 _0919_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_46_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1683_ _1683_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 _1683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1117_ _1136_/A _1121_/B vssd1 vssd1 vccd1 vccd1 _1119_/A sky130_fd_sc_hd__nand2_1
X_1048_ _1058_/B vssd1 vssd1 vccd1 vccd1 _1049_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1735_ _1735_/CLK _1735_/D vssd1 vssd1 vccd1 vccd1 _1735_/Q sky130_fd_sc_hd__dfxtp_1
X_1666_ _1666_/CLK _1666_/D vssd1 vssd1 vccd1 vccd1 _1666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627__65 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1697_/CLK sky130_fd_sc_hd__inv_2
X_1520_ hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1382_ _1588_/B _1382_/B vssd1 vssd1 vccd1 vccd1 _1383_/A sky130_fd_sc_hd__and2_1
X_1451_ _1451_/A hold88/A vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1718_ _1718_/CLK _1718_/D vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0951_ _1682_/Q _1670_/Q vssd1 vssd1 vccd1 vccd1 _0999_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0882_ _1682_/Q _1673_/Q vssd1 vssd1 vccd1 vccd1 _1358_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1503_ _1588_/B _1503_/B vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1296_ _1296_/A _1370_/C vssd1 vssd1 vccd1 vccd1 _1364_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1434_ _1434_/A hold56/A vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__nand2_1
X_1365_ _1301_/B _1361_/B _1364_/B vssd1 vssd1 vccd1 vccd1 _1370_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 rst vssd1 vssd1 vccd1 vccd1 _1700_/D sky130_fd_sc_hd__clkbuf_1
X_1150_ _1150_/A _1197_/A _1150_/C vssd1 vssd1 vccd1 vccd1 _1151_/C sky130_fd_sc_hd__nand3_1
X_1081_ _1353_/B vssd1 vssd1 vccd1 vccd1 _1082_/C sky130_fd_sc_hd__inv_2
X_0865_ _0865_/A vssd1 vssd1 vccd1 vccd1 _0866_/B sky130_fd_sc_hd__inv_2
X_0934_ _0995_/B _0935_/A _0985_/B vssd1 vssd1 vccd1 vccd1 _0982_/A sky130_fd_sc_hd__nand3_1
X_1417_ _1417_/A _1588_/B _1417_/C vssd1 vssd1 vccd1 vccd1 _1418_/A sky130_fd_sc_hd__and3_1
X_1348_ _1351_/A _1588_/B vssd1 vssd1 vccd1 vccd1 _1348_/Y sky130_fd_sc_hd__nand2_1
X_1279_ _1280_/B _1280_/A vssd1 vssd1 vccd1 vccd1 _1284_/A sky130_fd_sc_hd__or2_1
XFILLER_0_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1202_ _1246_/B vssd1 vssd1 vccd1 vccd1 _1203_/B sky130_fd_sc_hd__inv_2
X_1133_ _1133_/A _1197_/B vssd1 vssd1 vccd1 vccd1 _1137_/B sky130_fd_sc_hd__nand2_1
X_1064_ _1064_/A _1064_/B vssd1 vssd1 vccd1 vccd1 _1067_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0917_ _1141_/C _1141_/D _1163_/A _1163_/B vssd1 vssd1 vccd1 vccd1 _1079_/C sky130_fd_sc_hd__or4_1
X_0848_ _0849_/B _0849_/A vssd1 vssd1 vccd1 vccd1 _1293_/A sky130_fd_sc_hd__or2_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1682_ _1682_/CLK _1682_/D vssd1 vssd1 vccd1 vccd1 _1682_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1047_ _1055_/A _1056_/A vssd1 vssd1 vccd1 vccd1 _1058_/B sky130_fd_sc_hd__nand2_1
X_1116_ _1116_/A _1116_/B _1116_/C vssd1 vssd1 vccd1 vccd1 _1121_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_43_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1734_ _1734_/CLK _1734_/D vssd1 vssd1 vccd1 vccd1 _1734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1642__25 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1712_/CLK sky130_fd_sc_hd__inv_2
X_1450_ _1447_/X hold25/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__a21oi_1
X_1381_ _1381_/A vssd1 vssd1 vccd1 vccd1 _1718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1579_ _1579_/A hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1717_ _1717_/CLK _1717_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0950_ _1678_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _0999_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0881_ _1681_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__nand2_1
X_1502_ _1592_/A hold17/X vssd1 vssd1 vccd1 vccd1 _1685_/D sky130_fd_sc_hd__nor2_1
X_1433_ hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__inv_2
XFILLER_0_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1295_ _1294_/B _1295_/B _1295_/C vssd1 vssd1 vccd1 vccd1 _1370_/C sky130_fd_sc_hd__nand3b_2
X_1364_ _1361_/B _1364_/B _1364_/C vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ _1080_/A _1083_/A vssd1 vssd1 vccd1 vccd1 _1353_/B sky130_fd_sc_hd__nand2_1
X_0864_ _0864_/A vssd1 vssd1 vccd1 vccd1 _0866_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0933_ _0933_/A _0933_/B vssd1 vssd1 vccd1 vccd1 _0935_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1611__50 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1682_/CLK sky130_fd_sc_hd__inv_2
X_1416_ _1416_/A _1416_/B vssd1 vssd1 vccd1 vccd1 _1417_/C sky130_fd_sc_hd__nand2_1
X_1347_ _1347_/A _1347_/B vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__nand2_1
X_1278_ _1293_/A _1293_/B _1277_/A vssd1 vssd1 vccd1 vccd1 _1280_/A sky130_fd_sc_hd__o21ai_1
X_1656__6 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1726_/CLK sky130_fd_sc_hd__inv_2
X_1201_ _1201_/A _1241_/A vssd1 vssd1 vccd1 vccd1 _1246_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1132_ _1132_/A _1132_/B vssd1 vssd1 vccd1 vccd1 _1197_/B sky130_fd_sc_hd__nand2_1
X_1063_ _1065_/A _1112_/C vssd1 vssd1 vccd1 vccd1 _1064_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0916_ _1672_/Q vssd1 vssd1 vccd1 vccd1 _1163_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0847_ _1260_/A _1263_/D _1230_/B vssd1 vssd1 vccd1 vccd1 _0849_/A sky130_fd_sc_hd__or3_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_1681_ _1681_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _1681_/Q sky130_fd_sc_hd__dfxtp_2
X_1046_ _1055_/A _1056_/A vssd1 vssd1 vccd1 vccd1 _1132_/B sky130_fd_sc_hd__nor2_1
X_1115_ _1115_/A _1115_/B vssd1 vssd1 vccd1 vccd1 _1136_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1648__31 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1718_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_43_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1733_ _1733_/CLK _1733_/D vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1029_ _1094_/B _1031_/B vssd1 vssd1 vccd1 vccd1 _1159_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1380_ _1588_/B _1666_/Q vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__and2_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1618__56 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1688_/CLK sky130_fd_sc_hd__inv_2
X_1716_ _1716_/CLK _1716_/D vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
X_1578_ hold38/X _1579_/A vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__or2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0880_ _0886_/A _0901_/A vssd1 vssd1 vccd1 vccd1 _0885_/A sky130_fd_sc_hd__nand2_1
X_1501_ hold72/X vssd1 vssd1 vccd1 vccd1 _1686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1432_ _1432_/A _1458_/A vssd1 vssd1 vccd1 vccd1 _1434_/A sky130_fd_sc_hd__nor2_1
X_1363_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1724_/D sky130_fd_sc_hd__inv_2
X_1294_ _1294_/A _1294_/B vssd1 vssd1 vccd1 vccd1 _1296_/A sky130_fd_sc_hd__nand2_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0932_/A _0932_/B vssd1 vssd1 vccd1 vccd1 _0933_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0863_ _0863_/A _0863_/B vssd1 vssd1 vccd1 vccd1 _0902_/A sky130_fd_sc_hd__nand2_1
X_1415_ _1416_/B _1416_/A vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__or2_1
X_1346_ _1346_/A vssd1 vssd1 vccd1 vccd1 _1729_/D sky130_fd_sc_hd__clkbuf_1
X_1277_ _1277_/A _1277_/B vssd1 vssd1 vccd1 vccd1 _1293_/B sky130_fd_sc_hd__nand2_1
X_1200_ _1200_/A _1200_/B vssd1 vssd1 vccd1 vccd1 _1241_/A sky130_fd_sc_hd__or2_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ _1131_/A _1131_/B vssd1 vssd1 vccd1 vccd1 _1133_/A sky130_fd_sc_hd__nand2_1
X_1062_ _1112_/B _1062_/B _1062_/C vssd1 vssd1 vccd1 vccd1 _1112_/C sky130_fd_sc_hd__nand3_2
X_0915_ _1671_/Q vssd1 vssd1 vccd1 vccd1 _1163_/A sky130_fd_sc_hd__inv_2
X_0846_ _0846_/A vssd1 vssd1 vccd1 vccd1 _1230_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _1376_/A _1375_/B _1376_/B vssd1 vssd1 vccd1 vccd1 _1329_/Y sky130_fd_sc_hd__nand3_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_1680_ _1680_/CLK _1680_/D vssd1 vssd1 vccd1 vccd1 _1680_/Q sky130_fd_sc_hd__dfxtp_4
X_1114_ _1116_/B vssd1 vssd1 vccd1 vccd1 _1115_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1045_ _1667_/Q _1682_/Q vssd1 vssd1 vccd1 vccd1 _1056_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1663__13 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1733_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1732_ _1732_/CLK _1732_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
X_1594_ _1613_/A vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__buf_1
X_1028_ _1028_/A _1028_/B vssd1 vssd1 vccd1 vccd1 _1031_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1633__16 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1703_/CLK sky130_fd_sc_hd__inv_2
X_1715_ _1715_/CLK _1715_/D vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1577_/A _1583_/B vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__nor2_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1500_ _1500_/A _1588_/B hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__and3_1
X_1293_ _1293_/A _1293_/B vssd1 vssd1 vccd1 vccd1 _1294_/B sky130_fd_sc_hd__xnor2_1
X_1431_ hold83/A _1431_/B vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1362_ _1236_/A _1236_/B _1361_/X vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0931_ _0932_/B _0932_/A vssd1 vssd1 vccd1 vccd1 _0933_/A sky130_fd_sc_hd__or2_1
X_0862_ _0907_/B _0862_/B vssd1 vssd1 vccd1 vccd1 _0863_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1414_ _1414_/A _1414_/B vssd1 vssd1 vccd1 vccd1 _1416_/A sky130_fd_sc_hd__nand2_1
X_1276_ _1276_/A _1276_/B vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1345_ _1345_/A _1345_/B _1588_/B vssd1 vssd1 vccd1 vccd1 _1346_/A sky130_fd_sc_hd__and3_1
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1602__41 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1673_/CLK sky130_fd_sc_hd__inv_2
X_1130_ _1229_/B vssd1 vssd1 vccd1 vccd1 _1220_/B sky130_fd_sc_hd__inv_2
X_1061_ _1137_/A _1061_/B vssd1 vssd1 vccd1 vccd1 _1065_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0845_ _1670_/Q _1678_/Q vssd1 vssd1 vccd1 vccd1 _0846_/A sky130_fd_sc_hd__nand2_1
X_0914_ _1679_/Q vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__inv_2
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1259_ _1259_/A _1258_/Y vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__or2b_1
X_1328_ _1328_/A vssd1 vssd1 vccd1 vccd1 _1376_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1113_ _1134_/A _1113_/B vssd1 vssd1 vccd1 vccd1 _1116_/B sky130_fd_sc_hd__nand2_1
X_1044_ _1668_/Q _1681_/Q vssd1 vssd1 vccd1 vccd1 _1055_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1639__22 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1709_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_19_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1731_ _1731_/CLK _1731_/D vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfxtp_1
X_1593_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1593_/X sky130_fd_sc_hd__buf_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1027_ _1153_/B _1027_/B vssd1 vssd1 vccd1 vccd1 _1028_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1714_ _1714_/CLK _1714_/D vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
X_1576_ hold52/X _1576_/B vssd1 vssd1 vccd1 vccd1 _1583_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1623__61 _1630__68/A vssd1 vssd1 vccd1 vccd1 _1693_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1430_ _1701_/Q vssd1 vssd1 vccd1 vccd1 _1431_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ _1295_/B _1295_/C vssd1 vssd1 vccd1 vccd1 _1294_/A sky130_fd_sc_hd__nand2_1
X_1361_ _1700_/Q _1361_/B vssd1 vssd1 vccd1 vccd1 _1361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1559_ _1577_/A _1563_/A hold95/X vssd1 vssd1 vccd1 vccd1 _1560_/C sky130_fd_sc_hd__o21ai_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0930_ _0930_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0932_/A sky130_fd_sc_hd__nand2_1
X_0861_ _0871_/B vssd1 vssd1 vccd1 vccd1 _0862_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1413_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1702_/D sky130_fd_sc_hd__clkbuf_1
X_1275_ _1276_/B _1276_/A vssd1 vssd1 vccd1 vccd1 _1277_/A sky130_fd_sc_hd__or2_1
X_1344_ _1003_/A _1004_/B _1003_/C vssd1 vssd1 vccd1 vccd1 _1345_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1060_ _1112_/B _1062_/B vssd1 vssd1 vccd1 vccd1 _1137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0913_ _1680_/Q vssd1 vssd1 vccd1 vccd1 _1141_/C sky130_fd_sc_hd__inv_2
X_0844_ _1677_/Q vssd1 vssd1 vccd1 vccd1 _1263_/D sky130_fd_sc_hd__inv_2
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1189_ _1190_/B _1190_/A vssd1 vssd1 vccd1 vccd1 _1191_/A sky130_fd_sc_hd__or2_1
X_1258_ _1258_/A _1258_/B vssd1 vssd1 vccd1 vccd1 _1258_/Y sky130_fd_sc_hd__nand2_1
X_1327_ _1327_/A _1327_/B vssd1 vssd1 vccd1 vccd1 _1328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__0138_ clkbuf_0__0138_/X vssd1 vssd1 vccd1 vccd1 _1650__33/A sky130_fd_sc_hd__clkbuf_16
X_1112_ _1137_/C _1112_/B _1112_/C vssd1 vssd1 vccd1 vccd1 _1113_/B sky130_fd_sc_hd__nand3_1
X_1043_ _1132_/A _1043_/B vssd1 vssd1 vccd1 vccd1 _1050_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ _1592_/A hold37/X vssd1 vssd1 vccd1 vccd1 _1666_/D sky130_fd_sc_hd__nor2_1
X_1730_ _1730_/CLK _1730_/D vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
X_1026_ _1026_/A _1026_/B vssd1 vssd1 vccd1 vccd1 _1153_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ _1713_/CLK _1713_/D vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1575_ hold54/X vssd1 vssd1 vccd1 vccd1 _1670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1009_ _1020_/A _1021_/A vssd1 vssd1 vccd1 vccd1 _1154_/A sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1609__48 _1611__50/A vssd1 vssd1 vccd1 vccd1 _1680_/CLK sky130_fd_sc_hd__inv_2
X_1659__9 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1729_/CLK sky130_fd_sc_hd__inv_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1360_ _1360_/A vssd1 vssd1 vccd1 vccd1 _1725_/D sky130_fd_sc_hd__clkbuf_1
X_1291_ _1291_/A _1291_/B vssd1 vssd1 vccd1 vccd1 _1295_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ hold95/X _1577_/A _1563_/A vssd1 vssd1 vccd1 vccd1 _1560_/A sky130_fd_sc_hd__or3_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ hold30/X _1422_/B _1487_/A vssd1 vssd1 vccd1 vccd1 _1489_/X sky130_fd_sc_hd__a21o_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0860_ _0868_/A _0869_/A vssd1 vssd1 vccd1 vccd1 _0871_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1412_ _1588_/B input1/X vssd1 vssd1 vccd1 vccd1 _1413_/A sky130_fd_sc_hd__and2_1
X_1343_ _1343_/A vssd1 vssd1 vccd1 vccd1 _1730_/D sky130_fd_sc_hd__clkbuf_1
X_1274_ _1274_/A _1274_/B vssd1 vssd1 vccd1 vccd1 _1276_/A sky130_fd_sc_hd__xor2_1
X_0989_ _0953_/Y _0989_/B vssd1 vssd1 vccd1 vccd1 _0991_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0912_ _0922_/A _0930_/A vssd1 vssd1 vccd1 vccd1 _0920_/A sky130_fd_sc_hd__nand2_1
X_0843_ _1669_/Q vssd1 vssd1 vccd1 vccd1 _1260_/A sky130_fd_sc_hd__inv_2
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1326_ _1326_/A _1326_/B vssd1 vssd1 vccd1 vccd1 _1327_/B sky130_fd_sc_hd__nand2_1
X_1188_ _1188_/A _1188_/B vssd1 vssd1 vccd1 vccd1 _1190_/A sky130_fd_sc_hd__nand2_1
X_1257_ _1258_/A _1258_/B vssd1 vssd1 vccd1 vccd1 _1259_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1111_ _1112_/B _1137_/C vssd1 vssd1 vccd1 vccd1 _1134_/A sky130_fd_sc_hd__or2_1
X_1042_ _1054_/B vssd1 vssd1 vccd1 vccd1 _1043_/B sky130_fd_sc_hd__inv_2
Xmax_cap1 _0946_/A vssd1 vssd1 vccd1 vccd1 _1065_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1309_ _1310_/B _1310_/A vssd1 vssd1 vccd1 vccd1 _1318_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1591_ _1548_/Y _1590_/Y _1588_/B hold3/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
X_1025_ _1025_/A vssd1 vssd1 vccd1 vccd1 _1026_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1712_ _1712_/CLK _1712_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1574_ _1574_/A _1588_/B hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__and3_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1675_/Q _1674_/Q vssd1 vssd1 vccd1 vccd1 _1021_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1290_ _1290_/A vssd1 vssd1 vccd1 vccd1 _1291_/A sky130_fd_sc_hd__inv_2
X_1614__52 _1631__69/A vssd1 vssd1 vccd1 vccd1 _1684_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1557_ hold1/X hold13/X vssd1 vssd1 vccd1 vccd1 _1563_/A sky130_fd_sc_hd__nor2_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1486_/X hold34/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__a21oi_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1273_ _1273_/A _1273_/B vssd1 vssd1 vccd1 vccd1 _1274_/B sky130_fd_sc_hd__nor2_1
X_1411_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1703_/D sky130_fd_sc_hd__clkbuf_1
X_1342_ _1342_/A _1588_/B _1342_/C vssd1 vssd1 vccd1 vccd1 _1343_/A sky130_fd_sc_hd__and3_1
X_0988_ _0988_/A vssd1 vssd1 vccd1 vccd1 _1000_/A sky130_fd_sc_hd__inv_2
XFILLER_0_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0842_ _1274_/A _0842_/B vssd1 vssd1 vccd1 vccd1 _0849_/B sky130_fd_sc_hd__nand2_1
X_0911_ _0911_/A _0911_/B _0911_/C vssd1 vssd1 vccd1 vccd1 _0930_/A sky130_fd_sc_hd__or3_2
X_1256_ _1303_/A _1263_/D _0841_/B vssd1 vssd1 vccd1 vccd1 _1258_/B sky130_fd_sc_hd__or3b_1
X_1325_ _1376_/C vssd1 vssd1 vccd1 vccd1 _1375_/B sky130_fd_sc_hd__inv_2
X_1187_ _1187_/A _1671_/Q _1675_/Q vssd1 vssd1 vccd1 vccd1 _1190_/B sky130_fd_sc_hd__and3_1
XFILLER_0_37_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1110_ _1110_/A _1134_/B vssd1 vssd1 vccd1 vccd1 _1137_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1041_ _1051_/A _1052_/A vssd1 vssd1 vccd1 vccd1 _1054_/B sky130_fd_sc_hd__nand2_1
Xmax_cap2 _0940_/A vssd1 vssd1 vccd1 vccd1 _1034_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1239_ _1239_/A _1239_/B _1239_/C vssd1 vssd1 vccd1 vccd1 _1248_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1308_ _1318_/B _1307_/Y _1273_/A _1258_/Y _1259_/A vssd1 vssd1 vccd1 vccd1 _1310_/B
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_34_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1645__28 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1715_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1590_ hold73/X _1590_/B vssd1 vssd1 vccd1 vccd1 _1590_/Y sky130_fd_sc_hd__nor2_1
X_1024_ _1024_/A vssd1 vssd1 vccd1 vccd1 _1026_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__0138_ _1632_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__0138_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1711_ _1711_/CLK _1711_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1576_/B hold52/X _1585_/B vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__nand3_1
X_1007_ _1676_/Q _1673_/Q vssd1 vssd1 vccd1 vccd1 _1020_/A sky130_fd_sc_hd__nand2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1556_ hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__inv_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1487_/A hold33/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__nand2_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1651__1 _1659__9/A vssd1 vssd1 vccd1 vccd1 _1721_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1410_ _1588_/B input2/X vssd1 vssd1 vccd1 vccd1 _1411_/A sky130_fd_sc_hd__and2_1
XFILLER_0_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1272_ _1272_/A vssd1 vssd1 vccd1 vccd1 _1280_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1341_ _1341_/A _1341_/B vssd1 vssd1 vccd1 vccd1 _1342_/A sky130_fd_sc_hd__or2_1
XFILLER_0_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0987_ _0995_/A _0995_/B vssd1 vssd1 vccd1 vccd1 _0993_/A sky130_fd_sc_hd__nand2_1
X_1539_ hold43/X vssd1 vssd1 vccd1 vccd1 _1677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0841_ _0841_/A _0841_/B vssd1 vssd1 vccd1 vccd1 _0842_/B sky130_fd_sc_hd__nand2_1
X_0910_ _0926_/A _0910_/B vssd1 vssd1 vccd1 vccd1 _0922_/A sky130_fd_sc_hd__nand2_1
X_1186_ _1252_/B _1214_/C vssd1 vssd1 vccd1 vccd1 _1233_/B sky130_fd_sc_hd__nand2_1
X_1255_ _1260_/A _1303_/D _0841_/A vssd1 vssd1 vccd1 vccd1 _1258_/A sky130_fd_sc_hd__or3b_1
X_1324_ _1324_/A _1330_/A vssd1 vssd1 vccd1 vccd1 _1376_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ _1051_/A _1052_/A vssd1 vssd1 vccd1 vccd1 _1132_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1238_ _1237_/Y _1207_/B _1210_/B vssd1 vssd1 vccd1 vccd1 _1245_/A sky130_fd_sc_hd__o21ai_1
X_1169_ _1172_/A _1193_/A vssd1 vssd1 vccd1 vccd1 _1170_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1307_ _1307_/A _1307_/B vssd1 vssd1 vccd1 vccd1 _1307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1023_ _1153_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1710_ _1710_/CLK _1710_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_1572_ _1576_/B _1585_/B hold52/X vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__a21o_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1006_ _1079_/B _1079_/C vssd1 vssd1 vccd1 vccd1 _1078_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1555_ _1553_/X hold14/X _1592_/A vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__a21oi_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ hold33/X _1487_/A vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__or2_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1340_ _1340_/A vssd1 vssd1 vccd1 vccd1 _1731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1271_ _1259_/X _1267_/Y _1270_/Y vssd1 vssd1 vccd1 vccd1 _1272_/A sky130_fd_sc_hd__o21ai_1
X_0986_ _0986_/A _0997_/B vssd1 vssd1 vccd1 vccd1 _0995_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1469_ hold82/A hold88/A vssd1 vssd1 vccd1 vccd1 _1471_/A sky130_fd_sc_hd__nand2_1
X_1538_ _1538_/A _1588_/B hold42/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__and3_1
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0840_ _0841_/A _0841_/B vssd1 vssd1 vccd1 vccd1 _1274_/A sky130_fd_sc_hd__or2_1
X_1323_ _1323_/A _1323_/B vssd1 vssd1 vccd1 vccd1 _1330_/A sky130_fd_sc_hd__or2_1
X_1185_ _1251_/A vssd1 vssd1 vccd1 vccd1 _1214_/C sky130_fd_sc_hd__inv_2
X_1254_ _1295_/C _1288_/C vssd1 vssd1 vccd1 vccd1 _1287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0969_ _1062_/C vssd1 vssd1 vccd1 vccd1 _1061_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1306_ _1307_/A _1307_/B vssd1 vssd1 vccd1 vccd1 _1318_/B sky130_fd_sc_hd__or2_1
X_1237_ _1237_/A vssd1 vssd1 vccd1 vccd1 _1237_/Y sky130_fd_sc_hd__inv_2
X_1168_ _1168_/A _1188_/A _1168_/C vssd1 vssd1 vccd1 vccd1 _1193_/A sky130_fd_sc_hd__nand3_2
X_1099_ _1158_/A _1103_/B vssd1 vssd1 vccd1 vccd1 _1101_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ _1022_/A _1022_/B vssd1 vssd1 vccd1 vccd1 _1153_/A sky130_fd_sc_hd__nand2_1
X_1636__19 _1644__27/A vssd1 vssd1 vccd1 vccd1 _1706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650__33 _1650__33/A vssd1 vssd1 vccd1 vccd1 _1720_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_22_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ _1571_/A hold67/A vssd1 vssd1 vccd1 vccd1 _1576_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _0935_/A _0985_/B _0933_/B vssd1 vssd1 vccd1 vccd1 _1079_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput30 _1690_/Q vssd1 vssd1 vccd1 vccd1 p[5] sky130_fd_sc_hd__buf_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1554_ hold2/X _1577_/A hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o21ai_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1485_/A hold88/A vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__nand2_1
.ends

