* NGSPICE file created from lovers_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

.subckt lovers_controller becStatus[0] becStatus[1] becStatus[2] becStatus[3] data_in[0]
+ data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7]
+ data_in[8] data_in[9] data_out[0] data_out[10] data_out[11] data_out[12] data_out[13]
+ data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[1]
+ data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26]
+ data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] io_oeb io_out
+ ki la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6] la_data_in[7]
+ la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3]
+ la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ load_data load_status[0] load_status[1] load_status[2] load_status[3] load_status[4]
+ load_status[5] next_key slv_done slv_enable vccd1 vssd1 wb_clk_i wb_rst_i
XFILLER_0_185_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09671_ hold1368/X _16381_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _09003_/A hold433/X vssd1 vssd1 vccd1 vccd1 _15933_/D sky130_fd_sc_hd__and2_1
XFILLER_0_94_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08553_ _12420_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _15900_/D sky130_fd_sc_hd__and2_1
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08484_ _15217_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09105_ hold2374/X _09106_/B _09104_/Y _12984_/A vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ hold219/X hold724/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 hold340/A vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold351 hold351/A vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 hold373/A vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold384 hold67/X vssd1 vssd1 vccd1 vccd1 input16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold395 hold395/A vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14833_/C1 sky130_fd_sc_hd__buf_4
Xfanout831 fanout841/X vssd1 vssd1 vccd1 vccd1 _14859_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout842 _07787_/Y vssd1 vssd1 vccd1 vccd1 fanout842/X sky130_fd_sc_hd__buf_8
X_09938_ hold1408/X _16470_/Q _10022_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__mux2_1
Xfanout853 _11791_/A vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__buf_4
Xfanout864 _07783_/Y vssd1 vssd1 vccd1 vccd1 _15215_/A sky130_fd_sc_hd__clkbuf_16
Xfanout875 hold883/X vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__buf_8
Xfanout886 _15195_/A vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__clkbuf_16
X_09869_ hold1663/X hold3491/X _10481_/S vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__mux2_1
Xfanout897 hold667/X vssd1 vssd1 vccd1 vccd1 _14850_/A sky130_fd_sc_hd__buf_8
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 _08418_/X vssd1 vssd1 vccd1 vccd1 _15839_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 hold1148/X vssd1 vssd1 vccd1 vccd1 hold1149/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ hold2195/X hold5158/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__mux2_1
Xhold1062 _14299_/X vssd1 vssd1 vccd1 vccd1 _17949_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1073 _16183_/Q vssd1 vssd1 vccd1 vccd1 hold1073/X sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ hold1130/X hold3023/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__mux2_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _17894_/Q vssd1 vssd1 vccd1 vccd1 hold1084/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _07834_/X vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ hold2994/X hold3880/X _13793_/S vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ hold920/X _14554_/A2 _14549_/X _15044_/A vssd1 vssd1 vccd1 vccd1 hold921/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _17078_/Q _11762_/B _11762_/C vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and3_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ hold5203/X _13883_/B _13500_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _11103_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__or2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15000_/A _14481_/B vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ hold915/X _17055_/Q _11789_/C vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ _17453_/CLK _16220_/D vssd1 vssd1 vccd1 vccd1 _16220_/Q sky130_fd_sc_hd__dfxtp_1
X_13432_ hold4383/X _13814_/B _13431_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10644_ hold3642/X _10548_/A _10643_/X vssd1 vssd1 vccd1 vccd1 _10644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _17487_/CLK _16151_/D vssd1 vssd1 vccd1 vccd1 _16151_/Q sky130_fd_sc_hd__dfxtp_1
X_13363_ hold5130/X _13859_/B _13362_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13363_/X
+ sky130_fd_sc_hd__o211a_1
X_10575_ hold3673/X _11082_/A _10574_/X vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ hold5975/X _15109_/B hold541/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 hold542/A
+ sky130_fd_sc_hd__o211a_1
X_12314_ _12314_/A _12314_/B _12356_/C vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and3_1
XFILLER_0_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16082_ _17313_/CLK _16082_/D vssd1 vssd1 vccd1 vccd1 hold633/A sky130_fd_sc_hd__dfxtp_1
X_13294_ _13294_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ _15195_/A _18302_/Q hold302/X vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__mux2_1
X_12245_ hold1948/X hold4723/X _12341_/C vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ hold1712/X hold3372/X _12377_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11694_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__or2_1
X_16984_ _17896_/CLK _16984_/D vssd1 vssd1 vccd1 vccd1 _16984_/Q sky130_fd_sc_hd__dfxtp_1
X_15935_ _17345_/CLK _15935_/D vssd1 vssd1 vccd1 vccd1 hold611/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _11136_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17513_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10009_ _11203_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__nor2_1
X_15866_ _17649_/CLK _15866_/D vssd1 vssd1 vccd1 vccd1 _15866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14817_ hold1629/X _14828_/B _14816_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14817_/X
+ sky130_fd_sc_hd__o211a_1
X_17605_ _17701_/CLK _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _17731_/CLK _15797_/D vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17536_ _18380_/CLK _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14748_ _14980_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ _17482_/CLK _17467_/D vssd1 vssd1 vccd1 vccd1 _17467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14679_ hold2157/X _14666_/B _14678_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14679_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16418_ _18389_/CLK _16418_/D vssd1 vssd1 vccd1 vccd1 _16418_/Q sky130_fd_sc_hd__dfxtp_1
X_17398_ _18450_/CLK _17398_/D vssd1 vssd1 vccd1 vccd1 _17398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ _18360_/CLK _16349_/D vssd1 vssd1 vccd1 vccd1 _16349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6007 _18424_/Q vssd1 vssd1 vccd1 vccd1 hold6007/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6018 _09443_/Y vssd1 vssd1 vccd1 vccd1 _16307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold6029 la_data_in[21] vssd1 vssd1 vccd1 vccd1 hold570/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5306 _16328_/Q vssd1 vssd1 vccd1 vccd1 _13094_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_124_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5317 _10018_/Y vssd1 vssd1 vccd1 vccd1 _16496_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5328 _09535_/X vssd1 vssd1 vccd1 vccd1 _16335_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5339 _09526_/X vssd1 vssd1 vccd1 vccd1 _16332_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18019_ _18052_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4605 _16749_/Q vssd1 vssd1 vccd1 vccd1 hold4605/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4616 _11539_/X vssd1 vssd1 vccd1 vccd1 _17003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4627 _17060_/Q vssd1 vssd1 vccd1 vccd1 hold4627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4638 _11905_/X vssd1 vssd1 vccd1 vccd1 _17125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3904 _13846_/Y vssd1 vssd1 vccd1 vccd1 _17735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4649 _17025_/Q vssd1 vssd1 vccd1 vccd1 hold4649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3915 _16821_/Q vssd1 vssd1 vccd1 vccd1 hold3915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3926 _16352_/Q vssd1 vssd1 vccd1 vccd1 _13286_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3937 _10330_/X vssd1 vssd1 vccd1 vccd1 _16600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3948 _16814_/Q vssd1 vssd1 vccd1 vccd1 hold3948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3959 hold5872/X vssd1 vssd1 vccd1 vccd1 hold5873/A sky130_fd_sc_hd__buf_6
Xfanout149 _12836_/S vssd1 vssd1 vccd1 vccd1 _12800_/S sky130_fd_sc_hd__buf_4
X_07984_ _15553_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07984_/X sky130_fd_sc_hd__or2_1
X_09723_ _09918_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__or2_1
X_09654_ _09954_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__or2_1
X_08605_ hold35/X hold548/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08606_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09585_ _10491_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ hold407/X hold640/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__mux2_1
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ hold1225/X _08488_/B _08466_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ hold1010/X _08440_/A2 _08397_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10360_ hold4182/X _10589_/B _10359_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10360_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5840 _18405_/Q vssd1 vssd1 vccd1 vccd1 hold5840/X sky130_fd_sc_hd__dlygate4sd3_1
X_09019_ _12426_/A _09019_/B vssd1 vssd1 vccd1 vccd1 _16126_/D sky130_fd_sc_hd__and2_1
X_10291_ hold4609/X _10073_/B _10290_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10291_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5851 hold5851/A vssd1 vssd1 vccd1 vccd1 hold5851/X sky130_fd_sc_hd__clkbuf_4
Xhold5862 hold5944/X vssd1 vssd1 vccd1 vccd1 hold5862/X sky130_fd_sc_hd__buf_2
X_12030_ _12267_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__or2_1
Xhold5873 hold5873/A vssd1 vssd1 vccd1 vccd1 hold5873/X sky130_fd_sc_hd__clkbuf_4
Xhold5884 _07797_/X vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 la_data_in[19] vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5895 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold5895/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold192 hold295/X vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout650 _12927_/A vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_5_16__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_16__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
Xfanout661 _13627_/C1 vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__buf_4
Xfanout672 _08137_/A vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__buf_4
Xfanout683 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14171_/C1 sky130_fd_sc_hd__clkbuf_4
X_13981_ hold2127/X _13986_/B _13980_/Y _14350_/A vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout694 _08585_/A vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__buf_2
X_15720_ _17221_/CLK _15720_/D vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ hold3592/X _12931_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__mux2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _17878_/CLK _15651_/D vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ hold3331/X _12862_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _15103_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__or2_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18415_/CLK hold854/X vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__dfxtp_1
X_11814_ _12210_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__or2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _17282_/CLK _15582_/D vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ hold3528/X _12793_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__mux2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17321_ _17323_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _17321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _15105_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ hold3790/X _12093_/A _11744_/X vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _17252_/CLK _17252_/D vssd1 vssd1 vccd1 vccd1 _17252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464_ hold1195/X _14481_/B _14463_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14464_/X
+ sky130_fd_sc_hd__o211a_1
X_11676_ _12051_/A _11676_/B vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _17435_/CLK _16203_/D vssd1 vssd1 vccd1 vccd1 _16203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13415_ hold1010/X hold3217/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13416_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10627_ _11194_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/Y sky130_fd_sc_hd__nor2_1
X_17183_ _17282_/CLK _17183_/D vssd1 vssd1 vccd1 vccd1 _17183_/Q sky130_fd_sc_hd__dfxtp_1
X_14395_ _15129_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _18417_/CLK _16134_/D vssd1 vssd1 vccd1 vccd1 _16134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ hold1210/X hold3651/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__mux2_1
X_10558_ hold5170/X _10558_/A2 _10557_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _16676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16065_ _18413_/CLK _16065_/D vssd1 vssd1 vccd1 vccd1 hold716/A sky130_fd_sc_hd__dfxtp_1
X_13277_ _13276_/X hold3684/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__mux2_1
X_10489_ hold4743/X _10628_/B _10488_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10489_/X
+ sky130_fd_sc_hd__o211a_1
X_15016_ _15123_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15016_/X sky130_fd_sc_hd__or2_1
X_12228_ _12285_/A _12228_/B vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__or2_1
X_12159_ _12255_/A _12159_/B vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__or2_1
Xhold1809 _18093_/Q vssd1 vssd1 vccd1 vccd1 hold1809/X sky130_fd_sc_hd__dlygate4sd3_1
X_16967_ _17880_/CLK _16967_/D vssd1 vssd1 vccd1 vccd1 _16967_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _17513_/CLK _15918_/D vssd1 vssd1 vccd1 vccd1 hold553/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16898_ _18032_/CLK _16898_/D vssd1 vssd1 vccd1 vccd1 _16898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15849_ _17734_/CLK _15849_/D vssd1 vssd1 vccd1 vccd1 _15849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_266_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17584_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09370_ hold611/X _09367_/A _15447_/B1 hold707/X vssd1 vssd1 vccd1 vccd1 _09370_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ _15545_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08321_/Y sky130_fd_sc_hd__nand2_1
X_17519_ _17522_/CLK _17519_/D vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ _14866_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _14511_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5103 _13690_/X vssd1 vssd1 vccd1 vccd1 _17683_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5114 _16587_/Q vssd1 vssd1 vccd1 vccd1 hold5114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5125 _13594_/X vssd1 vssd1 vccd1 vccd1 _17651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5136 _17650_/Q vssd1 vssd1 vccd1 vccd1 hold5136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4402 _11635_/X vssd1 vssd1 vccd1 vccd1 _17035_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5147 _13492_/X vssd1 vssd1 vccd1 vccd1 _17617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4413 _16628_/Q vssd1 vssd1 vccd1 vccd1 hold4413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5158 _17124_/Q vssd1 vssd1 vccd1 vccd1 hold5158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5169 _13381_/X vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4424 _11884_/X vssd1 vssd1 vccd1 vccd1 _17118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4435 _16627_/Q vssd1 vssd1 vccd1 vccd1 hold4435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3701 _10648_/Y vssd1 vssd1 vccd1 vccd1 _16706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4446 _11980_/X vssd1 vssd1 vccd1 vccd1 _17150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3712 _09820_/X vssd1 vssd1 vccd1 vccd1 _16430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4457 _17189_/Q vssd1 vssd1 vccd1 vccd1 hold4457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3723 _10044_/Y vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4468 _09673_/X vssd1 vssd1 vccd1 vccd1 _16381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3734 _16541_/Q vssd1 vssd1 vccd1 vccd1 hold3734/X sky130_fd_sc_hd__buf_1
Xhold4479 _16688_/Q vssd1 vssd1 vccd1 vccd1 hold4479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3745 _16538_/Q vssd1 vssd1 vccd1 vccd1 hold3745/X sky130_fd_sc_hd__buf_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3756 hold4864/X vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3767 _17123_/Q vssd1 vssd1 vccd1 vccd1 hold3767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3778 _16904_/Q vssd1 vssd1 vccd1 vccd1 hold3778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3789 _11725_/Y vssd1 vssd1 vccd1 vccd1 _17065_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07967_ hold1457/X _07978_/B _07966_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _07967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ hold4319/X _10780_/A2 _09705_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__o211a_1
X_07898_ _15521_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07898_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09637_ hold5439/X _10025_/B _09636_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09637_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ hold5120/X _10070_/B _09567_/X _15144_/C1 vssd1 vssd1 vccd1 vccd1 _09568_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ _17523_/Q _17522_/Q vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__nor2_1
X_09499_ _18461_/Q _12510_/B vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_182_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11530_ hold3433/X _11617_/A2 _11529_/X _12666_/A vssd1 vssd1 vccd1 vccd1 _11530_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ hold4429/X _11747_/B _11460_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13193_/X _13199_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17543_/D sky130_fd_sc_hd__o21a_1
X_10412_ hold1489/X _16628_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11392_ hold4001/X _12338_/B _11391_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11392_/X
+ sky130_fd_sc_hd__o211a_1
X_14180_ _15199_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14180_/X sky130_fd_sc_hd__or2_1
X_13131_ _13130_/X hold3742/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__mux2_1
X_10343_ hold1344/X hold4129/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5670 _16502_/Q vssd1 vssd1 vccd1 vccd1 hold5670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5681 _16420_/Q vssd1 vssd1 vccd1 vccd1 hold5681/X sky130_fd_sc_hd__dlygate4sd3_1
X_10274_ hold1673/X hold4698/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__mux2_1
X_13062_ _13062_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__or2_1
Xhold5692 _10996_/X vssd1 vssd1 vccd1 vccd1 _16822_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12013_ hold4623/X _12299_/B _12012_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _12013_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4980 _10471_/X vssd1 vssd1 vccd1 vccd1 _16647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17870_ _17870_/CLK _17870_/D vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4991 _12073_/X vssd1 vssd1 vccd1 vccd1 _17181_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16821_ _18003_/CLK _16821_/D vssd1 vssd1 vccd1 vccd1 _16821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout480 _11219_/C vssd1 vssd1 vccd1 vccd1 _11789_/C sky130_fd_sc_hd__clkbuf_8
Xfanout491 _10763_/S vssd1 vssd1 vccd1 vccd1 _10874_/S sky130_fd_sc_hd__clkbuf_8
X_16752_ _18052_/CLK _16752_/D vssd1 vssd1 vccd1 vccd1 _16752_/Q sky130_fd_sc_hd__dfxtp_1
X_13964_ _15525_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13964_/X sky130_fd_sc_hd__or2_1
X_15703_ _17779_/CLK _15703_/D vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfxtp_1
X_12915_ _12918_/A _12915_/B vssd1 vssd1 vccd1 vccd1 _17481_/D sky130_fd_sc_hd__and2_1
X_16683_ _18268_/CLK _16683_/D vssd1 vssd1 vccd1 vccd1 _16683_/Q sky130_fd_sc_hd__dfxtp_1
X_13895_ _13897_/A _13895_/B vssd1 vssd1 vccd1 vccd1 _17755_/D sky130_fd_sc_hd__and2_1
XFILLER_0_158_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18422_ _18422_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _17275_/CLK _15634_/D vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12846_ _12849_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _17458_/D sky130_fd_sc_hd__and2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18353_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15565_ _17262_/CLK _15565_/D vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A _12777_/B vssd1 vssd1 vccd1 vccd1 _17435_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17318_/CLK _17304_/D vssd1 vssd1 vccd1 vccd1 hold398/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ hold2828/X _14554_/A2 _14515_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14516_/X
+ sky130_fd_sc_hd__o211a_1
X_18284_ _18378_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
X_11728_ _12301_/A _11728_/B vssd1 vssd1 vccd1 vccd1 _11728_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_154_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _15498_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__and2_1
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17235_ _17897_/CLK _17235_/D vssd1 vssd1 vccd1 vccd1 _17235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ hold607/X hold273/A vssd1 vssd1 vccd1 vccd1 _14447_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_153_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11659_ hold5344/X _11753_/B _11658_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17262_/CLK _17166_/D vssd1 vssd1 vccd1 vccd1 _17166_/Q sky130_fd_sc_hd__dfxtp_1
X_14378_ _14378_/A hold484/X vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold906 hold906/A vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16117_ _17340_/CLK _16117_/D vssd1 vssd1 vccd1 vccd1 hold676/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold917 hold917/A vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _13713_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__or2_1
Xhold928 hold928/A vssd1 vssd1 vccd1 vccd1 hold928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 hold939/A vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _17880_/CLK _17097_/D vssd1 vssd1 vccd1 vccd1 _17097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16048_ _16096_/CLK _16048_/D vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__dfxtp_1
Xhold3008 _17377_/Q vssd1 vssd1 vccd1 vccd1 hold3008/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3019 _12893_/X vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2307 _14717_/X vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08870_ hold23/X _16053_/Q _08932_/S vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__mux2_1
Xhold2318 _15584_/Q vssd1 vssd1 vccd1 vccd1 hold2318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 _13995_/X vssd1 vssd1 vccd1 vccd1 _17804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1606 _15652_/Q vssd1 vssd1 vccd1 vccd1 hold1606/X sky130_fd_sc_hd__dlygate4sd3_1
X_07821_ hold800/X _15551_/A _15553_/A vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__or3b_1
Xhold1617 hold6012/X vssd1 vssd1 vccd1 vccd1 _09472_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1628 _14153_/X vssd1 vssd1 vccd1 vccd1 _17880_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _18060_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1639 _08292_/X vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ _09438_/B _16297_/Q vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ _15547_/A hold335/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__or3_1
XFILLER_0_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ hold2830/X _08336_/A2 _08303_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _12804_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _16253_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ hold2820/X _08268_/B _08234_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08166_ _15517_/A hold1174/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ hold1968/X _08088_/B _08096_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _08097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4210 _10543_/X vssd1 vssd1 vccd1 vccd1 _16671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4221 _13354_/X vssd1 vssd1 vccd1 vccd1 _17571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4232 _16585_/Q vssd1 vssd1 vccd1 vccd1 hold4232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4243 _10240_/X vssd1 vssd1 vccd1 vccd1 _16570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4254 _16638_/Q vssd1 vssd1 vccd1 vccd1 hold4254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4265 hold5850/X vssd1 vssd1 vccd1 vccd1 hold5851/A sky130_fd_sc_hd__buf_4
Xhold3520 _17413_/Q vssd1 vssd1 vccd1 vccd1 hold3520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4276 _09754_/X vssd1 vssd1 vccd1 vccd1 _16408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3531 _16678_/Q vssd1 vssd1 vccd1 vccd1 hold3531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3542 _12764_/X vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4287 _16684_/Q vssd1 vssd1 vccd1 vccd1 hold4287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3553 _13486_/X vssd1 vssd1 vccd1 vccd1 _17615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4298 _10270_/X vssd1 vssd1 vccd1 vccd1 _16580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3564 _17713_/Q vssd1 vssd1 vccd1 vccd1 hold3564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2830 _15785_/Q vssd1 vssd1 vccd1 vccd1 hold2830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3575 _17363_/Q vssd1 vssd1 vccd1 vccd1 hold3575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 _16234_/Q vssd1 vssd1 vccd1 vccd1 hold2841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3586 _17356_/Q vssd1 vssd1 vccd1 vccd1 hold3586/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2852 _09093_/X vssd1 vssd1 vccd1 vccd1 _16161_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08999_ _13046_/C _08999_/B vssd1 vssd1 vccd1 vccd1 _09028_/S sky130_fd_sc_hd__or2_2
Xhold3597 _17355_/Q vssd1 vssd1 vccd1 vccd1 hold3597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2863 _14520_/X vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2874 _17755_/Q vssd1 vssd1 vccd1 vccd1 hold2874/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_188_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18080_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2885 _14597_/X vssd1 vssd1 vccd1 vccd1 _18092_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2896 _13953_/X vssd1 vssd1 vccd1 vccd1 _17783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_117_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18385_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ hold2660/X hold5548/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ hold1372/X _17411_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__mux2_1
X_13680_ _13770_/A _13680_/B vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ hold1488/X _16788_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__mux2_1
X_12631_ hold2481/X hold3014/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ hold523/X _09367_/A _15446_/B1 hold555/X vssd1 vssd1 vccd1 vccd1 _15350_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ hold2466/X _17365_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14301_ hold2801/X _14333_/A2 _14300_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14301_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11513_ hold773/X hold4941/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__mux2_1
X_15281_ _16292_/Q _15477_/A2 _15487_/B1 hold169/X _15280_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/D sky130_fd_sc_hd__a221o_1
X_12493_ hold56/X _12509_/A2 _12505_/A3 _12492_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold57/A sky130_fd_sc_hd__o311a_1
X_17020_ _17900_/CLK _17020_/D vssd1 vssd1 vccd1 vccd1 _17020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ _14913_/A hold273/X vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__nor2_1
X_11444_ hold1754/X hold3537/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14843_/A hold272/X vssd1 vssd1 vccd1 vccd1 _14206_/B sky130_fd_sc_hd__or2_4
X_11375_ hold2127/X _16949_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__mux2_1
X_13114_ _17565_/Q _17099_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__mux2_1
X_10326_ _10422_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__or2_1
X_14094_ _15547_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__nand2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _17524_/Q hold795/X _13044_/X _13056_/C _13048_/A vssd1 vssd1 vccd1 vccd1
+ hold796/A sky130_fd_sc_hd__o221a_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _18020_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_1
X_10257_ _10554_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10257_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _10380_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__or2_1
X_17853_ _17856_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
X_16804_ _18071_/CLK _16804_/D vssd1 vssd1 vccd1 vccd1 _16804_/Q sky130_fd_sc_hd__dfxtp_1
X_14996_ _15103_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__or2_1
X_17784_ _18432_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ _14627_/A hold273/A vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__or2_4
X_16735_ _18190_/CLK _16735_/D vssd1 vssd1 vccd1 vccd1 _16735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16666_ _18192_/CLK _16666_/D vssd1 vssd1 vccd1 vccd1 _16666_/Q sky130_fd_sc_hd__dfxtp_1
X_13878_ hold3931/X _13791_/A _13877_/X vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18405_ _18405_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
X_15617_ _17170_/CLK _15617_/D vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12829_ hold1994/X _17454_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__mux2_1
X_16597_ _18233_/CLK _16597_/D vssd1 vssd1 vccd1 vccd1 _16597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18336_ _18422_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ hold1857/X _15560_/A2 _15547_/Y _15502_/A vssd1 vssd1 vccd1 vccd1 _15548_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18267_ _18267_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _17323_/Q _15479_/A2 _09362_/C hold471/X _15478_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08020_ hold2681/X _08029_/B _08019_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _08020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17218_ _17703_/CLK _17218_/D vssd1 vssd1 vccd1 vccd1 _17218_/Q sky130_fd_sc_hd__dfxtp_1
X_18198_ _18198_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 hold714/A vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ _17744_/CLK _17149_/D vssd1 vssd1 vccd1 vccd1 _17149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold725 hold725/A vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/A vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__buf_12
Xhold758 hold758/A vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ hold978/X hold3463/X _10481_/S vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__mux2_1
Xhold769 hold779/X vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ hold65/X hold496/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2104 _17851_/Q vssd1 vssd1 vccd1 vccd1 hold2104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _18127_/Q vssd1 vssd1 vccd1 vccd1 hold2115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 _13985_/X vssd1 vssd1 vccd1 vccd1 _17799_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08853_ _12428_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _16045_/D sky130_fd_sc_hd__and2_1
Xhold2137 _15611_/Q vssd1 vssd1 vccd1 vccd1 hold2137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _18166_/Q vssd1 vssd1 vccd1 vccd1 hold1403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _14031_/X vssd1 vssd1 vccd1 vccd1 _17821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _18336_/Q vssd1 vssd1 vccd1 vccd1 hold2159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _15732_/Q vssd1 vssd1 vccd1 vccd1 hold1414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1425 _14518_/X vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 _18137_/Q vssd1 vssd1 vccd1 vccd1 hold1436/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_281_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18051_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__and2_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1447 _18069_/Q vssd1 vssd1 vccd1 vccd1 hold1447/X sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ _15473_/A hold106/X vssd1 vssd1 vccd1 vccd1 _16012_/D sky130_fd_sc_hd__and2_1
Xhold1458 _07967_/X vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _18174_/Q vssd1 vssd1 vccd1 vccd1 hold1469/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_210_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17903_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09405_ _07804_/A hold5895/X _15334_/A _09404_/X vssd1 vssd1 vccd1 vccd1 _09405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09336_ hold2656/X _09338_/A2 _09335_/X _12909_/A vssd1 vssd1 vccd1 vccd1 _09336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ hold235/X _16245_/Q _09277_/S vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08218_ hold1604/X _08213_/B _08217_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08218_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09198_ _15527_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _08149_/A _08149_/B vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11160_ hold3665/X _11640_/A _11159_/X vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__a21oi_1
Xhold4040 _10951_/X vssd1 vssd1 vccd1 vccd1 _16807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4051 _16629_/Q vssd1 vssd1 vccd1 vccd1 hold4051/X sky130_fd_sc_hd__dlygate4sd3_1
X_10111_ hold4349/X _10649_/B _10110_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10111_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4062 _10339_/X vssd1 vssd1 vccd1 vccd1 _16603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11091_ _11103_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11091_/X sky130_fd_sc_hd__or2_1
Xhold4073 _16597_/Q vssd1 vssd1 vccd1 vccd1 hold4073/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4084 _10129_/X vssd1 vssd1 vccd1 vccd1 _16533_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3350 _10150_/X vssd1 vssd1 vccd1 vccd1 _16540_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4095 _16699_/Q vssd1 vssd1 vccd1 vccd1 hold4095/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3361 _10141_/X vssd1 vssd1 vccd1 vccd1 _16537_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10042_ _11194_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/Y sky130_fd_sc_hd__nor2_1
Xhold3372 _17216_/Q vssd1 vssd1 vccd1 vccd1 hold3372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3383 _11239_/X vssd1 vssd1 vccd1 vccd1 _16903_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__buf_4
Xhold3394 _17072_/Q vssd1 vssd1 vccd1 vccd1 _11744_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2660 _18014_/Q vssd1 vssd1 vccd1 vccd1 hold2660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _14850_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__or2_1
Xhold2671 _13949_/X vssd1 vssd1 vccd1 vccd1 _17781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2682 _08020_/X vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2693 _18392_/Q vssd1 vssd1 vccd1 vccd1 hold2693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13801_ hold4032/X _13814_/B _13800_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _17720_/D
+ sky130_fd_sc_hd__o211a_1
Xhold1970 _18310_/Q vssd1 vssd1 vccd1 vccd1 hold1970/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ hold2149/X _14772_/B _14780_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14781_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1981 _15585_/Q vssd1 vssd1 vccd1 vccd1 hold1981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1992 _15790_/Q vssd1 vssd1 vccd1 vccd1 hold1992/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ hold1136/X _17155_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__mux2_1
X_16520_ _18205_/CLK _16520_/D vssd1 vssd1 vccd1 vccd1 _16520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ hold4055/X _13829_/B _13731_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13732_/X
+ sky130_fd_sc_hd__o211a_1
X_10944_ _11136_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__or2_1
X_16451_ _18388_/CLK _16451_/D vssd1 vssd1 vccd1 vccd1 _16451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13663_ hold5177/X _13883_/B _13662_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13663_/X
+ sky130_fd_sc_hd__o211a_1
X_10875_ _11106_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15402_ _15471_/A _15402_/B _15402_/C _15402_/D vssd1 vssd1 vccd1 vccd1 _15402_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_155_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12614_ hold3124/X _12613_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _18385_/CLK _16382_/D vssd1 vssd1 vccd1 vccd1 _16382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ hold5124/X _13880_/B _13593_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13594_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18217_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_85_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _15490_/A1 _15325_/X _15332_/X _15490_/B1 _18409_/Q vssd1 vssd1 vccd1 vccd1
+ _15333_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ hold3594/X _12544_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18052_ _18052_/CLK hold972/X vssd1 vssd1 vccd1 vccd1 hold971/A sky130_fd_sc_hd__dfxtp_1
X_15264_ _15334_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__and2_1
X_12476_ _17331_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__or2_1
X_17003_ _17884_/CLK _17003_/D vssd1 vssd1 vccd1 vccd1 _17003_/Q sky130_fd_sc_hd__dfxtp_1
X_14215_ hold2344/X _14198_/B _14214_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14215_/X
+ sky130_fd_sc_hd__o211a_1
X_11427_ _12018_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
XANTENNA_5 _13076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _15195_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _15545_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nand2_1
X_11358_ _11649_/A _11358_/B vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ hold4759/X _10619_/B _10308_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__o211a_1
X_14077_ hold773/X _14105_/A2 _14076_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 hold774/A
+ sky130_fd_sc_hd__o211a_1
X_11289_ _11694_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__or2_1
X_13028_ _13029_/B _13039_/A _13028_/C vssd1 vssd1 vccd1 vccd1 _13028_/X sky130_fd_sc_hd__and3b_1
X_17905_ _17905_/CLK hold844/X vssd1 vssd1 vccd1 vccd1 hold843/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _17887_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _17799_/CLK _17767_/D vssd1 vssd1 vccd1 vccd1 _17767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14979_ hold952/X _15006_/B _14978_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 hold953/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16718_ _18062_/CLK _16718_/D vssd1 vssd1 vccd1 vccd1 _16718_/Q sky130_fd_sc_hd__dfxtp_1
X_17698_ _17730_/CLK _17698_/D vssd1 vssd1 vccd1 vccd1 _17698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16649_ _18315_/CLK _16649_/D vssd1 vssd1 vccd1 vccd1 _16649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09121_ hold800/X _09121_/B _15553_/A _15551_/A vssd1 vssd1 vccd1 vccd1 hold801/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18319_ _18319_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ hold65/X hold477/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ _14511_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold511 hold511/A vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold533 hold533/A vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 hold544/A vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 hold555/A vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 hold566/A vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 hold577/A vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold588 hold588/A vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__or2_1
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _12428_/A _08905_/B vssd1 vssd1 vccd1 vccd1 _16070_/D sky130_fd_sc_hd__and2_1
X_09885_ _09981_/A _09885_/B vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__or2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _14480_/X vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _08459_/X vssd1 vssd1 vccd1 vccd1 _15858_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ hold214/X hold420/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08837_/B sky130_fd_sc_hd__mux2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _15720_/Q vssd1 vssd1 vccd1 vccd1 hold1222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _18202_/Q vssd1 vssd1 vccd1 vccd1 hold1233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 _18063_/Q vssd1 vssd1 vccd1 vccd1 hold1244/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1255 _18271_/Q vssd1 vssd1 vccd1 vccd1 hold1255/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 _14079_/X vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _18320_/Q vssd1 vssd1 vccd1 vccd1 hold1277/X sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ hold219/X hold720/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__mux2_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _17833_/Q vssd1 vssd1 vccd1 vccd1 hold1288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _15188_/X vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _12438_/A _08698_/B vssd1 vssd1 vccd1 vccd1 _15970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ hold4822/X _11732_/B _10659_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _10660_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _15541_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10591_ _10651_/A _10591_/B vssd1 vssd1 vccd1 vccd1 _10591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ hold5239/X _12234_/A _12329_/X vssd1 vssd1 vccd1 vccd1 _12330_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12261_ _12267_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _14681_/A hold272/X vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__nor2_1
X_11212_ _12331_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12192_ _13797_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11143_ _11155_/A _11143_/B vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__nor2_1
Xoutput75 _13153_/A vssd1 vssd1 vccd1 vccd1 output75/X sky130_fd_sc_hd__buf_6
XFILLER_0_128_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput86 _13233_/A vssd1 vssd1 vccd1 vccd1 output86/X sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_132_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18382_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput97 _13081_/A vssd1 vssd1 vccd1 vccd1 output97/X sky130_fd_sc_hd__buf_6
X_15951_ _16128_/CLK _15951_/D vssd1 vssd1 vccd1 vccd1 hold699/A sky130_fd_sc_hd__dfxtp_1
X_11074_ _11168_/A _11735_/B _11073_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _11074_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3180 _10602_/Y vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10025_ _16499_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__and3_1
Xhold3191 _17115_/Q vssd1 vssd1 vccd1 vccd1 hold3191/X sky130_fd_sc_hd__dlygate4sd3_1
X_14902_ _14972_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__or2_1
X_15882_ _17592_/CLK _15882_/D vssd1 vssd1 vccd1 vccd1 _15882_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2490 _17982_/Q vssd1 vssd1 vccd1 vccd1 hold2490/X sky130_fd_sc_hd__dlygate4sd3_1
X_17621_ _17749_/CLK _17621_/D vssd1 vssd1 vccd1 vccd1 _17621_/Q sky130_fd_sc_hd__dfxtp_1
X_14833_ hold1688/X _14828_/B _14832_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _18223_/CLK _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _15103_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14764_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _13392_/A _11976_/B vssd1 vssd1 vccd1 vccd1 _11976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _18360_/CLK _16503_/D vssd1 vssd1 vccd1 vccd1 _16503_/Q sky130_fd_sc_hd__dfxtp_1
X_13715_ hold2725/X hold4959/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__mux2_1
X_17483_ _17484_/CLK _17483_/D vssd1 vssd1 vccd1 vccd1 _17483_/Q sky130_fd_sc_hd__dfxtp_1
X_10927_ hold5668/X _11213_/B _10926_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10927_/X
+ sky130_fd_sc_hd__o211a_1
X_14695_ hold2959/X _14720_/B _14694_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16434_ _18373_/CLK _16434_/D vssd1 vssd1 vccd1 vccd1 _16434_/Q sky130_fd_sc_hd__dfxtp_1
X_13646_ hold1227/X _17669_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13647_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10858_ hold4494/X _11726_/B _10857_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _10858_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _18420_/CLK _16365_/D vssd1 vssd1 vccd1 vccd1 _16365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ hold1638/X _17646_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13578_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10789_ hold3275/X _11747_/B _10788_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10789_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15316_ _17335_/Q _15486_/B1 _15485_/B1 hold350/X vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__a22o_1
X_18104_ _18220_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
X_12528_ _12936_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _17352_/D sky130_fd_sc_hd__and2_1
XFILLER_0_48_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16296_ _16314_/CLK _16296_/D vssd1 vssd1 vccd1 vccd1 _16296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15247_ hold391/X _09357_/A _15484_/B1 hold393/X _15246_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18035_ _18035_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ hold26/X _12445_/A _12505_/A3 _12458_/X _12420_/A vssd1 vssd1 vccd1 vccd1
+ hold27/A sky130_fd_sc_hd__o311a_1
Xhold4809 _17257_/Q vssd1 vssd1 vccd1 vccd1 hold4809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15178_ hold2818/X _15161_/B _15177_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15178_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ hold5961/X _14148_/B _14128_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14129_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout309 fanout337/X vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__clkbuf_4
X_09670_ hold3287/X _10070_/B _09669_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ hold136/X hold432/X _08655_/S vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__mux2_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17819_ _17884_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08552_ hold53/X hold524/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ hold2006/X _08488_/B _08482_/Y _08373_/A vssd1 vssd1 vccd1 vccd1 _08483_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _15219_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _15414_/A hold413/X vssd1 vssd1 vccd1 vccd1 _16134_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 data_in[14] vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 hold352/A vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold374 hold374/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 input16/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold396 hold396/A vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _15144_/C1 vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout821 _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14867_/C1 sky130_fd_sc_hd__buf_4
X_09937_ hold5502/X _10049_/B _09936_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09937_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout832 _14955_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_5_15__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
Xfanout843 _13864_/A vssd1 vssd1 vccd1 vccd1 _13822_/A sky130_fd_sc_hd__buf_8
Xfanout854 _10651_/A vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__buf_6
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout865 _15109_/A vssd1 vssd1 vccd1 vccd1 _15543_/A sky130_fd_sc_hd__buf_12
Xfanout876 hold883/X vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__clkbuf_16
Xfanout887 hold1157/X vssd1 vssd1 vccd1 vccd1 hold1158/A sky130_fd_sc_hd__buf_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09868_ hold5588/X _10780_/A2 _09867_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09868_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout898 _14972_/A vssd1 vssd1 vccd1 vccd1 _15513_/A sky130_fd_sc_hd__buf_8
Xhold1030 hold1071/X vssd1 vssd1 vccd1 vccd1 hold1030/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _15791_/Q vssd1 vssd1 vccd1 vccd1 hold1041/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08819_ _15244_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _16028_/D sky130_fd_sc_hd__and2_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 hold1150/X vssd1 vssd1 vccd1 vccd1 hold1052/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 _18362_/Q vssd1 vssd1 vccd1 vccd1 hold1063/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ hold3855/X _10028_/B _09798_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09799_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 _09141_/X vssd1 vssd1 vccd1 vccd1 _16183_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _14183_/X vssd1 vssd1 vccd1 vccd1 _17894_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 hold1259/X vssd1 vssd1 vccd1 vccd1 hold1260/A sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ hold3267/X _12308_/B _11829_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _12343_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__nor2_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13788_/A _13500_/B vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__or2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ hold1704/X hold3708/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__mux2_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ hold1199/X _14481_/B _14479_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14480_/X
+ sky130_fd_sc_hd__o211a_1
X_11692_ hold5506/X _12329_/B _11691_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11692_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13431_ _13800_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__or2_1
X_10643_ _16705_/Q _10643_/B _10643_/C vssd1 vssd1 vccd1 vccd1 _10643_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ _17487_/CLK _16150_/D vssd1 vssd1 vccd1 vccd1 _16150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _13764_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ _10574_/A _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__and3_1
X_15101_ hold540/X _15125_/B vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__or2_1
XFILLER_0_133_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12313_ _13822_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12313_/Y sky130_fd_sc_hd__nor2_1
X_16081_ _18405_/CLK _16081_/D vssd1 vssd1 vccd1 vccd1 hold482/A sky130_fd_sc_hd__dfxtp_1
X_13293_ _13292_/X hold3642/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15032_ _15032_/A _15032_/B vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_313_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17692_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12244_ _12338_/A _12347_/B _12243_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _12244_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12175_ hold4490/X _13844_/B _12174_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12175_/X
+ sky130_fd_sc_hd__o211a_1
X_11126_ hold1447/X hold5662/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__mux2_1
X_16983_ _17895_/CLK _16983_/D vssd1 vssd1 vccd1 vccd1 _16983_/Q sky130_fd_sc_hd__dfxtp_1
X_15934_ _17524_/CLK _15934_/D vssd1 vssd1 vccd1 vccd1 hold726/A sky130_fd_sc_hd__dfxtp_1
X_11057_ hold2967/X hold5570/X _11153_/C vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10008_ _13134_/A _09924_/A _10007_/X vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__a21oi_1
X_15865_ _17703_/CLK _15865_/D vssd1 vssd1 vccd1 vccd1 _15865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17604_ _17739_/CLK _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14816_ _15209_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__or2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _17730_/CLK _15796_/D vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _18308_/CLK _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11959_ hold4818/X _12341_/B _11958_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11959_/X
+ sky130_fd_sc_hd__o211a_1
X_14747_ hold2897/X _14774_/B _14746_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17466_ _17484_/CLK _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/Q sky130_fd_sc_hd__dfxtp_1
X_14678_ _14786_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14678_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16417_ _18330_/CLK _16417_/D vssd1 vssd1 vccd1 vccd1 _16417_/Q sky130_fd_sc_hd__dfxtp_1
X_13629_ _13734_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17397_ _18450_/CLK _17397_/D vssd1 vssd1 vccd1 vccd1 _17397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6008 _18421_/Q vssd1 vssd1 vccd1 vccd1 hold6008/X sky130_fd_sc_hd__dlygate4sd3_1
X_16348_ _18315_/CLK _16348_/D vssd1 vssd1 vccd1 vccd1 _16348_/Q sky130_fd_sc_hd__dfxtp_1
Xhold6019 _16313_/Q vssd1 vssd1 vccd1 vccd1 hold6019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ _17485_/CLK _16279_/D vssd1 vssd1 vccd1 vccd1 _16279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5307 _09993_/Y vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5318 _16738_/Q vssd1 vssd1 vccd1 vccd1 hold5318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5329 _16771_/Q vssd1 vssd1 vccd1 vccd1 hold5329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4606 _10681_/X vssd1 vssd1 vccd1 vccd1 _16717_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18018_ _18052_/CLK hold772/X vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4617 _16938_/Q vssd1 vssd1 vccd1 vccd1 hold4617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4628 _11614_/X vssd1 vssd1 vccd1 vccd1 _17028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4639 _17176_/Q vssd1 vssd1 vccd1 vccd1 hold4639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3905 hold5834/X vssd1 vssd1 vccd1 vccd1 hold3905/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3916 _10897_/X vssd1 vssd1 vccd1 vccd1 _16789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3927 _10065_/Y vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3938 _16791_/Q vssd1 vssd1 vccd1 vccd1 hold3938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3949 _10876_/X vssd1 vssd1 vccd1 vccd1 _16782_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07983_ hold1548/X _07978_/B _07982_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ hold980/X hold3861/X _09893_/S vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09653_ hold2524/X hold3562/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__mux2_1
X_08604_ _15314_/A hold678/X vssd1 vssd1 vccd1 vccd1 _15924_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09584_ hold1580/X _13286_/A _10628_/C vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__mux2_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08535_ _15344_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _15891_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08466_ _15199_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08397_ hold892/X _08445_/B vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ hold443/X hold714/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5830 hold5830/A vssd1 vssd1 vccd1 vccd1 hold5830/X sky130_fd_sc_hd__buf_2
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ _10506_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/X sky130_fd_sc_hd__or2_1
Xhold5841 hold5841/A vssd1 vssd1 vccd1 vccd1 hold5841/X sky130_fd_sc_hd__buf_2
Xhold5852 _16283_/Q vssd1 vssd1 vccd1 vccd1 hold5852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5863 hold5863/A vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_12
XFILLER_0_131_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5874 hold5947/X vssd1 vssd1 vccd1 vccd1 hold5874/X sky130_fd_sc_hd__buf_2
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5885 hold6035/X vssd1 vssd1 vccd1 vccd1 _09447_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 input47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5896 _16905_/Q vssd1 vssd1 vccd1 vccd1 hold5896/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold297/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__buf_4
Xfanout640 fanout660/X vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__buf_2
Xfanout651 _12927_/A vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__buf_4
Xfanout662 _13627_/C1 vssd1 vssd1 vccd1 vccd1 _13801_/C1 sky130_fd_sc_hd__clkbuf_4
X_13980_ _15000_/A _13980_/B vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__nand2_1
Xfanout673 _08137_/A vssd1 vssd1 vccd1 vccd1 _13411_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout684 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__buf_4
XFILLER_0_77_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout695 _12984_/A vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__buf_4
X_12931_ hold2628/X hold3042/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12931_/X sky130_fd_sc_hd__mux2_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _18445_/CLK _15650_/D vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfxtp_1
X_12862_ hold2462/X hold3289/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11813_ hold1222/X hold3165/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__mux2_1
X_14601_ hold1696/X _14612_/B _14600_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14601_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _17217_/CLK _15581_/D vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ hold2605/X hold3119/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__mux2_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _18421_/CLK hold33/X vssd1 vssd1 vccd1 vccd1 _17320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ hold2394/X _14554_/A2 _14531_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _14532_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11744_/A _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__and3_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17251_ _17283_/CLK _17251_/D vssd1 vssd1 vccd1 vccd1 _17251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14463_ _14517_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14463_/X sky130_fd_sc_hd__or2_1
X_11675_ hold1320/X hold5381/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ hold4161/X _13814_/B _13413_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13414_/X
+ sky130_fd_sc_hd__o211a_1
X_16202_ _17435_/CLK _16202_/D vssd1 vssd1 vccd1 vccd1 _16202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10626_ hold3639/X _10548_/A _10625_/X vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__a21oi_1
X_17182_ _17584_/CLK _17182_/D vssd1 vssd1 vccd1 vccd1 _17182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14394_ hold207/X hold273/A vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__or2_4
XFILLER_0_181_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ _18408_/CLK _16133_/D vssd1 vssd1 vccd1 vccd1 hold391/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13345_ hold3336/X _13832_/B _13344_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _18407_/CLK _16064_/D vssd1 vssd1 vccd1 vccd1 hold555/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13276_ hold5266/X _13275_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__mux2_2
X_10488_ _10491_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10488_/X sky130_fd_sc_hd__or2_1
X_15015_ hold2232/X _15006_/B _15014_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ hold1008/X _17233_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ hold1273/X _17210_/Q _13388_/S vssd1 vssd1 vccd1 vccd1 _12159_/B sky130_fd_sc_hd__mux2_1
X_11109_ _11115_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__or2_1
X_12089_ hold1954/X _17187_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__mux2_1
X_16966_ _17878_/CLK _16966_/D vssd1 vssd1 vccd1 vccd1 _16966_/Q sky130_fd_sc_hd__dfxtp_1
X_15917_ _18408_/CLK _15917_/D vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16897_ _18070_/CLK _16897_/D vssd1 vssd1 vccd1 vccd1 _16897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _17734_/CLK hold742/X vssd1 vssd1 vccd1 vccd1 _15848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15779_ _17678_/CLK _15779_/D vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ hold1877/X _08323_/B _08319_/Y _12756_/A vssd1 vssd1 vccd1 vccd1 _08320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ _17522_/CLK hold903/X vssd1 vssd1 vccd1 vccd1 _17518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ hold2082/X _08262_/B _08250_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08251_/X
+ sky130_fd_sc_hd__o211a_1
X_17449_ _17456_/CLK _17449_/D vssd1 vssd1 vccd1 vccd1 _17449_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_235_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17281_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08182_ hold1634/X _08209_/B _08181_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5104 _17714_/Q vssd1 vssd1 vccd1 vccd1 hold5104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5115 _10195_/X vssd1 vssd1 vccd1 vccd1 _16555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5126 _17238_/Q vssd1 vssd1 vccd1 vccd1 hold5126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5137 _13495_/X vssd1 vssd1 vccd1 vccd1 _17618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4403 _16960_/Q vssd1 vssd1 vccd1 vccd1 hold4403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5148 _16550_/Q vssd1 vssd1 vccd1 vccd1 hold5148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4414 _10318_/X vssd1 vssd1 vccd1 vccd1 _16596_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5159 _11806_/X vssd1 vssd1 vccd1 vccd1 _17092_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4425 _16970_/Q vssd1 vssd1 vccd1 vccd1 hold4425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4436 _10315_/X vssd1 vssd1 vccd1 vccd1 _16595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4447 _17094_/Q vssd1 vssd1 vccd1 vccd1 hold4447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3702 _16910_/Q vssd1 vssd1 vccd1 vccd1 hold3702/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4458 _12001_/X vssd1 vssd1 vccd1 vccd1 _17157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3713 _16928_/Q vssd1 vssd1 vccd1 vccd1 hold3713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3724 _10045_/Y vssd1 vssd1 vccd1 vccd1 _16505_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4469 _17008_/Q vssd1 vssd1 vccd1 vccd1 hold4469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3735 _10632_/Y vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3746 _10623_/Y vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3757 _10596_/Y vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3768 _12378_/Y vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3779 _11721_/Y vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07966_ _08311_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09705_ _10779_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__or2_1
X_07897_ hold2650/X _07918_/B _07896_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _07897_/X
+ sky130_fd_sc_hd__o211a_1
X_09636_ _09924_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _09975_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08518_ hold1828/X _08503_/Y _08517_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _08518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09498_ _14681_/A _09498_/B _09498_/C _09498_/D vssd1 vssd1 vccd1 vccd1 _12510_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ _08504_/A _14913_/A vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__or2_4
XFILLER_0_68_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11460_ _11652_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ hold4510/X _10619_/B _10410_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11391_ _12051_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__or2_1
X_13130_ _17567_/Q _17101_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ hold4518/X _10589_/B _10341_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10342_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5660 _11104_/X vssd1 vssd1 vccd1 vccd1 _16858_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13061_ _13060_/X hold5170/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
X_10273_ hold4779/X _10628_/B _10272_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _10273_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5671 _09940_/X vssd1 vssd1 vccd1 vccd1 _16470_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5682 _09694_/X vssd1 vssd1 vccd1 vccd1 _16388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5693 _17046_/Q vssd1 vssd1 vccd1 vccd1 hold5693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12012_ _12204_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4970 _13666_/X vssd1 vssd1 vccd1 vccd1 _17675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4981 _17243_/Q vssd1 vssd1 vccd1 vccd1 hold4981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4992 _16969_/Q vssd1 vssd1 vccd1 vccd1 hold4992/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_39_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18305_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16820_ _18055_/CLK _16820_/D vssd1 vssd1 vccd1 vccd1 _16820_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout470 fanout484/X vssd1 vssd1 vccd1 vccd1 _12368_/C sky130_fd_sc_hd__buf_4
Xfanout481 _11219_/C vssd1 vssd1 vccd1 vccd1 _11765_/C sky130_fd_sc_hd__clkbuf_8
Xfanout492 _09893_/S vssd1 vssd1 vccd1 vccd1 _10010_/C sky130_fd_sc_hd__clkbuf_8
X_16751_ _18020_/CLK _16751_/D vssd1 vssd1 vccd1 vccd1 _16751_/Q sky130_fd_sc_hd__dfxtp_1
X_13963_ hold1235/X _13980_/B _13962_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _13963_/X
+ sky130_fd_sc_hd__o211a_1
X_15702_ _17898_/CLK _15702_/D vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ hold3270/X _12913_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__mux2_1
X_13894_ _14218_/A hold2874/X hold244/X vssd1 vssd1 vccd1 vccd1 _13895_/B sky130_fd_sc_hd__mux2_1
X_16682_ _18353_/CLK _16682_/D vssd1 vssd1 vccd1 vccd1 _16682_/Q sky130_fd_sc_hd__dfxtp_1
X_18421_ _18421_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
X_15633_ _17253_/CLK _15633_/D vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfxtp_1
X_12845_ hold3063/X _12844_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__mux2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18388_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ hold3455/X _12775_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__mux2_1
X_15564_ _17232_/CLK _15564_/D vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17318_/CLK _17303_/D vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11727_ hold3719/X _11631_/A _11726_/X vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14515_ _14980_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14515_/X sky130_fd_sc_hd__or2_1
X_18283_ _18315_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ hold892/X hold1034/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _17902_/CLK _17234_/D vssd1 vssd1 vccd1 vccd1 _17234_/Q sky130_fd_sc_hd__dfxtp_1
X_11658_ _11658_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11658_/X sky130_fd_sc_hd__or2_1
X_14446_ hold2036/X hold209/X _14445_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10609_ _10651_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _10609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _17252_/CLK _17165_/D vssd1 vssd1 vccd1 vccd1 _17165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14377_ hold335/X hold483/X hold275/X vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__mux2_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11589_ _12036_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold907 hold907/A vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ _17343_/CLK _16116_/D vssd1 vssd1 vccd1 vccd1 hold534/A sky130_fd_sc_hd__dfxtp_1
X_13328_ hold1838/X hold3150/X _13808_/C vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__mux2_1
Xhold918 hold918/A vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17096_ _17128_/CLK _17096_/D vssd1 vssd1 vccd1 vccd1 _17096_/Q sky130_fd_sc_hd__dfxtp_1
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_16047_ _18308_/CLK _16047_/D vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__dfxtp_1
X_13259_ _13258_/X _16925_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__mux2_1
Xhold3009 _12602_/X vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2308 _17932_/Q vssd1 vssd1 vccd1 vccd1 hold2308/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2319 _07878_/X vssd1 vssd1 vccd1 vccd1 _15584_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07820_ hold270/X _14555_/C _14735_/A _09495_/C vssd1 vssd1 vccd1 vccd1 _09122_/A
+ sky130_fd_sc_hd__or4_1
Xhold1607 _08022_/X vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _18054_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1618 _09425_/X vssd1 vssd1 vccd1 vccd1 _16298_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 _18198_/Q vssd1 vssd1 vccd1 vccd1 hold1629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16949_ _17829_/CLK _16949_/D vssd1 vssd1 vccd1 vccd1 _16949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _07804_/A _09463_/B _15304_/A _09420_/X vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09352_ hold86/X hold265/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09366_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_75_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08303_ _15527_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ _15559_/A hold2120/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08234_ _14740_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ _08355_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _14728_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__or2_1
Xhold4200 _17580_/Q vssd1 vssd1 vccd1 vccd1 hold4200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4211 _16769_/Q vssd1 vssd1 vccd1 vccd1 hold4211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4222 _16570_/Q vssd1 vssd1 vccd1 vccd1 hold4222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4233 _10189_/X vssd1 vssd1 vccd1 vccd1 _16553_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4244 _16973_/Q vssd1 vssd1 vccd1 vccd1 hold4244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3510 _12244_/X vssd1 vssd1 vccd1 vccd1 _17238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4255 _10348_/X vssd1 vssd1 vccd1 vccd1 _16606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4266 _09388_/X vssd1 vssd1 vccd1 vccd1 _16282_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3521 _17147_/Q vssd1 vssd1 vccd1 vccd1 hold3521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4277 _17024_/Q vssd1 vssd1 vccd1 vccd1 hold4277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3532 _10468_/X vssd1 vssd1 vccd1 vccd1 _16646_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3543 _16677_/Q vssd1 vssd1 vccd1 vccd1 hold3543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4288 _10486_/X vssd1 vssd1 vccd1 vccd1 _16652_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4299 _16660_/Q vssd1 vssd1 vccd1 vccd1 hold4299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3554 _16646_/Q vssd1 vssd1 vccd1 vccd1 hold3554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2820 _15752_/Q vssd1 vssd1 vccd1 vccd1 hold2820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3565 _13684_/X vssd1 vssd1 vccd1 vccd1 _17681_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2831 _08304_/X vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3576 _12560_/X vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08998_ _09003_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _16116_/D sky130_fd_sc_hd__and2_1
Xhold2842 _15756_/Q vssd1 vssd1 vccd1 vccd1 hold2842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3587 _17491_/Q vssd1 vssd1 vccd1 vccd1 hold3587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3598 _16331_/Q vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2853 _17976_/Q vssd1 vssd1 vccd1 vccd1 hold2853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 _17400_/Q vssd1 vssd1 vccd1 vccd1 hold2864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2875 _18203_/Q vssd1 vssd1 vccd1 vccd1 hold2875/X sky130_fd_sc_hd__dlygate4sd3_1
X_07949_ hold1214/X _07991_/A2 _07948_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _07949_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2886 _17757_/Q vssd1 vssd1 vccd1 vccd1 hold2886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2897 _18164_/Q vssd1 vssd1 vccd1 vccd1 hold2897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ hold3940/X _11150_/B _10959_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__o211a_1
X_09619_ hold3999/X _10001_/B _09618_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__o211a_1
X_10891_ hold4250/X _11177_/B _10890_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12630_ _12855_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _17386_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_157_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _12933_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _17363_/D sky130_fd_sc_hd__and2_1
XFILLER_0_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ hold4647/X _11792_/B _11511_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11512_/X
+ sky130_fd_sc_hd__o211a_1
X_14300_ _14980_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14300_/X sky130_fd_sc_hd__or2_1
X_15280_ hold216/X _15486_/A2 _15446_/B1 _16057_/Q vssd1 vssd1 vccd1 vccd1 _15280_/X
+ sky130_fd_sc_hd__a22o_1
X_12492_ _17339_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ hold1872/X _14216_/Y _14230_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11443_ hold4745/X _11732_/B _11442_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ _14843_/A hold272/X vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__nor2_1
X_11374_ hold5409/X _11762_/B _11373_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _11374_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ _13113_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__and2_1
X_10325_ hold2293/X hold3219/X _10523_/S vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__mux2_1
X_14093_ hold2104/X _14094_/B _14092_/Y _14356_/A vssd1 vssd1 vccd1 vccd1 _14093_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _17518_/Q hold927/X _13043_/X _13030_/A vssd1 vssd1 vccd1 vccd1 _13044_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5490 _16746_/Q vssd1 vssd1 vccd1 vccd1 hold5490/X sky130_fd_sc_hd__dlygate4sd3_1
X_17921_ _18062_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_1
X_10256_ hold1515/X hold4359/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__mux2_1
X_17852_ _17852_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
X_10187_ hold1723/X hold4093/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__mux2_1
X_16803_ _18070_/CLK _16803_/D vssd1 vssd1 vccd1 vccd1 _16803_/Q sky130_fd_sc_hd__dfxtp_1
X_17783_ _18432_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
X_14995_ hold1698/X _15006_/B _14994_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _14995_/X
+ sky130_fd_sc_hd__o211a_1
X_16734_ _18025_/CLK _16734_/D vssd1 vssd1 vccd1 vccd1 _16734_/Q sky130_fd_sc_hd__dfxtp_1
X_13946_ _14627_/A hold273/A vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__nor2_2
X_16665_ _18095_/CLK _16665_/D vssd1 vssd1 vccd1 vccd1 _16665_/Q sky130_fd_sc_hd__dfxtp_1
X_13877_ _17746_/Q _13880_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__and3_1
XFILLER_0_158_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _18421_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _17584_/CLK _15616_/D vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _12843_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _17452_/D sky130_fd_sc_hd__and2_1
X_16596_ _18218_/CLK _16596_/D vssd1 vssd1 vccd1 vccd1 _16596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18335_ _18337_/CLK hold542/X vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15547_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12759_ _12813_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _17429_/D sky130_fd_sc_hd__and2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ _18266_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
X_15478_ hold432/X _09367_/A _09392_/C hold565/X vssd1 vssd1 vccd1 vccd1 _15478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _17217_/CLK _17217_/D vssd1 vssd1 vccd1 vccd1 _17217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14429_ _15543_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14429_/Y sky130_fd_sc_hd__nand2_1
X_18197_ _18197_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 hold704/A vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ _17584_/CLK _17148_/D vssd1 vssd1 vccd1 vccd1 _17148_/Q sky130_fd_sc_hd__dfxtp_1
Xhold715 hold715/A vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold726 hold726/A vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 hold737/A vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ hold5183/X _10628_/B _09969_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09970_/X
+ sky130_fd_sc_hd__o211a_1
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _17895_/CLK _17079_/D vssd1 vssd1 vccd1 vccd1 _17079_/Q sky130_fd_sc_hd__dfxtp_1
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ _15304_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _16078_/D sky130_fd_sc_hd__and2_1
XFILLER_0_21_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2105 _14093_/X vssd1 vssd1 vccd1 vccd1 _17851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2116 _14669_/X vssd1 vssd1 vccd1 vccd1 _18127_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08852_ hold251/X hold328/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__mux2_1
Xhold2127 _17797_/Q vssd1 vssd1 vccd1 vccd1 hold2127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2138 _07935_/X vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _18181_/Q vssd1 vssd1 vccd1 vccd1 hold2149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 _14751_/X vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _08192_/X vssd1 vssd1 vccd1 vccd1 _15732_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07803_ _07804_/B _07801_/B _07802_/Y vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__o21ai_1
Xhold1426 _15731_/Q vssd1 vssd1 vccd1 vccd1 hold1426/X sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ hold65/X _16012_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__mux2_1
Xhold1437 _14691_/X vssd1 vssd1 vccd1 vccd1 _18137_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1448 _14546_/X vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _16269_/Q vssd1 vssd1 vccd1 vccd1 hold1459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _09438_/B _09404_/B vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_250_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _15557_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09266_ _09272_/A hold115/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08217_ _14330_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09197_ hold2605/X _09218_/B _09196_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _09197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08148_ _14726_/A hold1848/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ hold2189/X _08088_/B _08078_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _08079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4030 _16603_/Q vssd1 vssd1 vccd1 vccd1 hold4030/X sky130_fd_sc_hd__dlygate4sd3_1
X_10110_ _10554_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__or2_1
Xhold4041 _17585_/Q vssd1 vssd1 vccd1 vccd1 hold4041/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4052 _10321_/X vssd1 vssd1 vccd1 vccd1 _16597_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4063 _16406_/Q vssd1 vssd1 vccd1 vccd1 hold4063/X sky130_fd_sc_hd__dlygate4sd3_1
X_11090_ hold2713/X _16854_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _11091_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4074 _10225_/X vssd1 vssd1 vccd1 vccd1 _16565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3340 _17191_/Q vssd1 vssd1 vccd1 vccd1 hold3340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4085 _16705_/Q vssd1 vssd1 vccd1 vccd1 hold4085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4096 _10531_/X vssd1 vssd1 vccd1 vccd1 _16667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3351 _17061_/Q vssd1 vssd1 vccd1 vccd1 hold3351/X sky130_fd_sc_hd__dlygate4sd3_1
X_10041_ _13222_/A _10380_/A _10040_/X vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3362 _17144_/Q vssd1 vssd1 vccd1 vccd1 hold3362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3373 _16881_/Q vssd1 vssd1 vccd1 vccd1 hold3373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__buf_2
Xhold3384 _17412_/Q vssd1 vssd1 vccd1 vccd1 hold3384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2650 _15592_/Q vssd1 vssd1 vccd1 vccd1 hold2650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3395 _11650_/X vssd1 vssd1 vccd1 vccd1 _17040_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__clkbuf_4
Xhold2661 _14432_/X vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 _18359_/Q vssd1 vssd1 vccd1 vccd1 hold2672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2683 _18090_/Q vssd1 vssd1 vccd1 vccd1 hold2683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__buf_1
Xhold2694 _15220_/X vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1960 _15581_/Q vssd1 vssd1 vccd1 vccd1 hold1960/X sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _13800_/A _13800_/B vssd1 vssd1 vccd1 vccd1 _13800_/X sky130_fd_sc_hd__or2_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__buf_4
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _15227_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__or2_1
X_11992_ hold4945/X _13844_/B _11991_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11992_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1971 _15801_/Q vssd1 vssd1 vccd1 vccd1 hold1971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1982 _07880_/X vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1993 _08314_/X vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13731_ _13734_/A _13731_/B vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__or2_1
X_10943_ hold2822/X _16805_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__mux2_1
X_16450_ _18395_/CLK _16450_/D vssd1 vssd1 vccd1 vccd1 _16450_/Q sky130_fd_sc_hd__dfxtp_1
X_13662_ _13788_/A _13662_/B vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10874_ hold911/X _16782_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__mux2_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _16304_/Q _09362_/A _09392_/B hold552/X _15400_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_38_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _18433_/Q hold3037/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__mux2_1
X_16381_ _18390_/CLK _16381_/D vssd1 vssd1 vccd1 vccd1 _16381_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13593_ _13791_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13593_/X sky130_fd_sc_hd__or2_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18126_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_1
X_15332_ _15489_/A _15332_/B _15332_/C _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/X
+ sky130_fd_sc_hd__or4_1
X_12544_ hold1646/X hold3236/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ _18051_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12475_ hold71/X _12509_/A2 _12505_/A3 _12474_/X _15374_/A vssd1 vssd1 vccd1 vccd1
+ hold72/A sky130_fd_sc_hd__o311a_1
X_15263_ _15490_/A1 _15255_/X _15262_/X _15490_/B1 hold3844/X vssd1 vssd1 vccd1 vccd1
+ _15263_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _17882_/CLK _17002_/D vssd1 vssd1 vccd1 vccd1 _17002_/Q sky130_fd_sc_hd__dfxtp_1
X_14214_ _15559_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__or2_1
X_11426_ hold1201/X hold4629/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15194_ hold3010/X _15221_/B _15193_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14145_ hold1818/X _14148_/B _14144_/Y _13905_/A vssd1 vssd1 vccd1 vccd1 _14145_/X
+ sky130_fd_sc_hd__o211a_1
X_11357_ hold1889/X _16943_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11358_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10308_ _10524_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__or2_1
X_14076_ hold747/X _14106_/B vssd1 vssd1 vccd1 vccd1 _14076_/X sky130_fd_sc_hd__or2_1
X_11288_ hold1683/X hold5356/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__mux2_1
X_13027_ _13034_/D hold901/X vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__and2_1
X_17904_ _17904_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_1
X_10239_ _10554_/A _10239_/B vssd1 vssd1 vccd1 vccd1 _10239_/X sky130_fd_sc_hd__or2_1
X_17835_ _17855_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
X_17766_ _18064_/CLK _17766_/D vssd1 vssd1 vccd1 vccd1 _17766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14978_ hold826/X _15018_/B vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717_ _17984_/CLK _16717_/D vssd1 vssd1 vccd1 vccd1 _16717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _13929_/A hold282/X vssd1 vssd1 vccd1 vccd1 _17772_/D sky130_fd_sc_hd__and2_1
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17697_ _17697_/CLK _17697_/D vssd1 vssd1 vccd1 vccd1 _17697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16648_ _18214_/CLK _16648_/D vssd1 vssd1 vccd1 vccd1 _16648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16579_ _18230_/CLK _16579_/D vssd1 vssd1 vccd1 vccd1 _16579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09120_ _18459_/Q _11155_/A _18462_/Q vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nor3_1
X_18318_ _18382_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09051_ _15344_/A _09051_/B vssd1 vssd1 vccd1 vccd1 _16142_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _18383_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08002_ hold1654/X _08033_/B _08001_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _08002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold501 data_in[12] vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold512 hold512/A vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold523 hold523/A vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold534 hold534/A vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 hold545/A vssd1 vssd1 vccd1 vccd1 input14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 hold556/A vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold567 hold567/A vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 hold578/A vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ hold987/X hold4549/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__mux2_1
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_14__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_90_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ hold184/X hold461/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08905_/B sky130_fd_sc_hd__mux2_1
X_09884_ hold2098/X _16452_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _17814_/Q vssd1 vssd1 vccd1 vccd1 hold1201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _18148_/Q vssd1 vssd1 vccd1 vccd1 hold1212/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _12438_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _16036_/D sky130_fd_sc_hd__and2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _18454_/Q vssd1 vssd1 vccd1 vccd1 hold1223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 _14825_/X vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 _14534_/X vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1256 _14971_/X vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _18364_/Q vssd1 vssd1 vccd1 vccd1 hold1267/X sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ _15344_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _16003_/D sky130_fd_sc_hd__and2_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1278 _15646_/Q vssd1 vssd1 vccd1 vccd1 hold1278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 _14057_/X vssd1 vssd1 vccd1 vccd1 _17833_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08697_ hold214/X hold392/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08698_/B sky130_fd_sc_hd__mux2_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ hold1459/X _09325_/B _09317_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _09318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ hold3693/X _10551_/A _10589_/X vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09249_ _15525_/A hold2541/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12260_ hold1269/X _17244_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_133_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ hold3601/X _11115_/A _11210_/X vssd1 vssd1 vccd1 vccd1 _11211_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ hold1832/X hold4184/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__mux2_1
X_11142_ hold3610/X _11061_/A _11141_/X vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput76 _13161_/A vssd1 vssd1 vccd1 vccd1 output76/X sky130_fd_sc_hd__buf_6
Xoutput87 _13241_/A vssd1 vssd1 vccd1 vccd1 output87/X sky130_fd_sc_hd__buf_6
X_15950_ _18425_/CLK _15950_/D vssd1 vssd1 vccd1 vccd1 hold649/A sky130_fd_sc_hd__dfxtp_1
X_11073_ _11640_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__or2_1
Xoutput98 _13089_/A vssd1 vssd1 vccd1 vccd1 output98/X sky130_fd_sc_hd__buf_6
Xhold3170 _12328_/Y vssd1 vssd1 vccd1 vccd1 _17266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3181 _10603_/Y vssd1 vssd1 vccd1 vccd1 _16691_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10024_ _11155_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _10024_/Y sky130_fd_sc_hd__nor2_1
X_14901_ hold1576/X hold657/X _14900_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _14901_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3192 _12354_/Y vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__dlygate4sd3_1
X_15881_ _17719_/CLK hold963/X vssd1 vssd1 vccd1 vccd1 hold962/A sky130_fd_sc_hd__dfxtp_1
X_17620_ _17748_/CLK _17620_/D vssd1 vssd1 vccd1 vccd1 _17620_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2480 _15703_/Q vssd1 vssd1 vccd1 vccd1 hold2480/X sky130_fd_sc_hd__dlygate4sd3_1
X_14832_ _15225_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14832_/X sky130_fd_sc_hd__or2_1
Xhold2491 _18005_/Q vssd1 vssd1 vccd1 vccd1 hold2491/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_172_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _18095_/CLK _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1790 _18039_/Q vssd1 vssd1 vccd1 vccd1 hold1790/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ hold1720/X _14774_/B _14762_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14763_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11975_ hold2143/X hold5106/X _13871_/C vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__mux2_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _18319_/CLK _16502_/D vssd1 vssd1 vccd1 vccd1 _16502_/Q sky130_fd_sc_hd__dfxtp_1
X_13714_ hold3402/X _13808_/B _13713_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _13714_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17482_ _17482_/CLK _17482_/D vssd1 vssd1 vccd1 vccd1 _17482_/Q sky130_fd_sc_hd__dfxtp_1
X_10926_ _11103_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__or2_1
X_14694_ _14980_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ _18378_/CLK _16433_/D vssd1 vssd1 vccd1 vccd1 _16433_/Q sky130_fd_sc_hd__dfxtp_1
X_13645_ hold4559/X _13856_/B _13644_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13645_/X
+ sky130_fd_sc_hd__o211a_1
X_10857_ _11631_/A _10857_/B vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16364_ _18334_/CLK _16364_/D vssd1 vssd1 vccd1 vccd1 _16364_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ hold3322/X _13862_/B _13575_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13576_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _11076_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18103_ _18231_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_1
X_15315_ hold308/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12527_ hold3436/X _12526_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16295_ _16314_/CLK _16295_/D vssd1 vssd1 vccd1 vccd1 _16295_/Q sky130_fd_sc_hd__dfxtp_1
X_18034_ _18034_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _17328_/Q _15486_/B1 _15485_/B1 hold329/X vssd1 vssd1 vccd1 vccd1 _15246_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _17322_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _11697_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__or2_1
X_12389_ hold32/X hold449/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__mux2_1
X_15177_ _15231_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14128_ hold883/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14059_ hold1079/X _14105_/A2 _14058_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14059_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ _09011_/A hold602/X vssd1 vssd1 vccd1 vccd1 _15932_/D sky130_fd_sc_hd__and2_1
X_17818_ _17884_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _12420_/A _08551_/B vssd1 vssd1 vccd1 vccd1 _15899_/D sky130_fd_sc_hd__and2_1
X_17749_ _17749_/CLK _17749_/D vssd1 vssd1 vccd1 vccd1 _17749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08482_ _15541_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ hold2048/X _09106_/B _09102_/Y _12987_/A vssd1 vssd1 vccd1 vccd1 _09103_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ hold184/X _16134_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold413/A sky130_fd_sc_hd__mux2_1
XFILLER_0_142_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 hold70/X vssd1 vssd1 vccd1 vccd1 input10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold487/X vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold375 hold375/A vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 hold386/A vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14941_/C1 sky130_fd_sc_hd__buf_4
Xhold397 hold397/A vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _15144_/C1 vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__buf_2
X_09936_ _09954_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__or2_1
Xfanout822 fanout841/X vssd1 vssd1 vccd1 vccd1 _14863_/C1 sky130_fd_sc_hd__buf_4
Xfanout833 _14955_/C1 vssd1 vssd1 vccd1 vccd1 _14869_/C1 sky130_fd_sc_hd__buf_4
Xfanout844 _13864_/A vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__buf_8
Xfanout855 _11791_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__buf_8
Xfanout866 _15109_/A vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__buf_8
Xfanout877 hold882/X vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__buf_6
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _11106_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09867_/X sky130_fd_sc_hd__or2_1
Xhold1020 _18082_/Q vssd1 vssd1 vccd1 vccd1 hold1020/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 hold826/X vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__buf_8
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1031 hold1031/A vssd1 vssd1 vccd1 vccd1 _15123_/A sky130_fd_sc_hd__buf_12
Xfanout899 _15187_/A vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__buf_8
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 _08316_/X vssd1 vssd1 vccd1 vccd1 _15791_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ hold47/X hold376/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__mux2_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 hold1053/A vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__buf_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 _15158_/X vssd1 vssd1 vccd1 vccd1 _18362_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _09918_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__or2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 _16149_/Q vssd1 vssd1 vccd1 vccd1 hold1075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _17971_/Q vssd1 vssd1 vccd1 vccd1 hold1086/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 hold1261/X vssd1 vssd1 vccd1 vccd1 hold1097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ hold443/X hold452/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__mux2_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ hold5365/X _11670_/A _11759_/X vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__a21oi_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ hold5340/X _11216_/B _10710_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10711_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ _12234_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__or2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10642_ _10651_/A _10642_/B vssd1 vssd1 vccd1 vccd1 _10642_/Y sky130_fd_sc_hd__nor2_1
X_13430_ hold2546/X _17597_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13361_ hold1280/X hold3793/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _11194_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10573_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15100_ hold2856/X _15109_/B _15099_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _15100_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12312_ hold3880/X _13794_/A _12311_/X vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__a21oi_1
X_16080_ _17331_/CLK _16080_/D vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
X_13292_ hold3705/X _13291_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13292_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__or2_1
X_15031_ _15193_/A hold3060/X hold302/X vssd1 vssd1 vccd1 vccd1 _15032_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ _13749_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11125_ hold5651/X _11222_/B _11124_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _11125_/X
+ sky130_fd_sc_hd__o211a_1
X_16982_ _17798_/CLK _16982_/D vssd1 vssd1 vccd1 vccd1 _16982_/Q sky130_fd_sc_hd__dfxtp_1
X_15933_ _17343_/CLK _15933_/D vssd1 vssd1 vccd1 vccd1 hold432/A sky130_fd_sc_hd__dfxtp_1
X_11056_ hold3961/X _11150_/B _11055_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__o211a_1
X_10007_ _16493_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__and3_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ _17735_/CLK hold909/X vssd1 vssd1 vccd1 vccd1 hold908/A sky130_fd_sc_hd__dfxtp_1
X_17603_ _17669_/CLK _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
X_14815_ hold2183/X _14822_/B _14814_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14815_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _17634_/CLK _15795_/D vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17534_ _18380_/CLK _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _15193_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14746_/X sky130_fd_sc_hd__or2_1
X_11958_ _12246_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17465_ _17484_/CLK _17465_/D vssd1 vssd1 vccd1 vccd1 _17465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10909_ hold5108/X _11177_/B _10908_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o211a_1
X_14677_ hold2141/X _14664_/B _14676_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__o211a_1
X_11889_ _12279_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16416_ _18330_/CLK _16416_/D vssd1 vssd1 vccd1 vccd1 _16416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ hold1934/X hold4067/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17396_ _18448_/CLK _17396_/D vssd1 vssd1 vccd1 vccd1 _17396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _18396_/CLK _16347_/D vssd1 vssd1 vccd1 vccd1 _16347_/Q sky130_fd_sc_hd__dfxtp_1
X_13559_ hold2369/X hold5066/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6009 _18417_/Q vssd1 vssd1 vccd1 vccd1 hold6009/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _17480_/CLK _16278_/D vssd1 vssd1 vccd1 vccd1 _16278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5308 _09994_/Y vssd1 vssd1 vccd1 vccd1 _16488_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5319 _11223_/Y vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__dlygate4sd3_1
X_18017_ _18337_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
X_15229_ _15229_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__or2_1
Xhold4607 _16439_/Q vssd1 vssd1 vccd1 vccd1 hold4607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4618 _11248_/X vssd1 vssd1 vccd1 vccd1 _16906_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4629 _16966_/Q vssd1 vssd1 vccd1 vccd1 hold4629/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3906 _15253_/X vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3917 _16397_/Q vssd1 vssd1 vccd1 vccd1 hold3917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3928 _10066_/Y vssd1 vssd1 vccd1 vccd1 _16512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3939 _10807_/X vssd1 vssd1 vccd1 vccd1 _16759_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07982_ _15551_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07982_/X sky130_fd_sc_hd__or2_1
X_09721_ hold5354/X _10025_/B _09720_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09721_/X
+ sky130_fd_sc_hd__o211a_1
X_09652_ hold4063/X _10571_/B _09651_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09652_/X
+ sky130_fd_sc_hd__o211a_1
X_08603_ hold407/X hold677/X _08661_/S vssd1 vssd1 vccd1 vccd1 hold678/A sky130_fd_sc_hd__mux2_1
X_09583_ hold5038/X _10073_/B _09582_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ hold68/X hold447/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08535_/B sky130_fd_sc_hd__mux2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ hold1128/X _08488_/B _08464_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ hold2431/X _08440_/A2 _08395_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09017_ _15454_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _16125_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5820 hold5897/X vssd1 vssd1 vccd1 vccd1 hold5820/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5831 _18400_/Q vssd1 vssd1 vccd1 vccd1 hold5831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5842 _18408_/Q vssd1 vssd1 vccd1 vccd1 hold5842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5853 hold5853/A vssd1 vssd1 vccd1 vccd1 hold5853/X sky130_fd_sc_hd__clkbuf_4
Xhold5864 _18418_/Q vssd1 vssd1 vccd1 vccd1 hold5864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5875 hold5875/A vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_12
Xhold161 hold52/X vssd1 vssd1 vccd1 vccd1 input6/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5886 _16322_/Q vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5897 _17518_/Q vssd1 vssd1 vccd1 vccd1 hold5897/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 input47/X vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold183 hold410/X vssd1 vssd1 vccd1 vccd1 hold411/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold280/X vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout630 _07824_/Y vssd1 vssd1 vccd1 vccd1 _15477_/A2 sky130_fd_sc_hd__buf_6
Xfanout641 _12810_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__clkbuf_4
X_09919_ hold5401/X _10013_/B _09918_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout652 _12927_/A vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__buf_2
Xfanout663 _13627_/C1 vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__buf_4
Xfanout674 fanout842/X vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__clkbuf_4
Xfanout685 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14510_/C1 sky130_fd_sc_hd__buf_4
Xfanout696 _12984_/A vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__buf_4
X_12930_ _12933_/A _12930_/B vssd1 vssd1 vccd1 vccd1 _17486_/D sky130_fd_sc_hd__and2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ _12924_/A _12861_/B vssd1 vssd1 vccd1 vccd1 _17463_/D sky130_fd_sc_hd__and2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _15209_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__or2_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ hold4311/X _12308_/B _11811_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11812_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _17283_/CLK _15580_/D vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12825_/A _12792_/B vssd1 vssd1 vccd1 vccd1 _17440_/D sky130_fd_sc_hd__and2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _15103_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__or2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _12301_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11743_/Y sky130_fd_sc_hd__nor2_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17282_/CLK _17250_/D vssd1 vssd1 vccd1 vccd1 _17250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ hold2971/X _14487_/B _14461_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14462_/X
+ sky130_fd_sc_hd__o211a_1
X_11674_ _11768_/A _11798_/B _11673_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11674_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ _17484_/CLK _16201_/D vssd1 vssd1 vccd1 vccd1 _16201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ _13800_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ _16699_/Q _10643_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__and3_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ _17744_/CLK _17181_/D vssd1 vssd1 vccd1 vccd1 _17181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14393_ hold207/X hold273/A vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16132_ _18417_/CLK _16132_/D vssd1 vssd1 vccd1 vccd1 _16132_/Q sky130_fd_sc_hd__dfxtp_1
X_13344_ _13737_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ hold2570/X hold5142/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _17329_/CLK _16063_/D vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__dfxtp_1
X_10487_ hold2415/X hold4196/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10488_/B sky130_fd_sc_hd__mux2_1
X_13275_ _13274_/X hold5321/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13275_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _15229_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__or2_1
X_12226_ hold4909/X _12311_/B _12225_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ hold5046/X _12347_/B _12156_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ hold1244/X _16860_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__mux2_1
X_12088_ hold4737/X _13844_/B _12087_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__o211a_1
X_16965_ _17877_/CLK _16965_/D vssd1 vssd1 vccd1 vccd1 _16965_/Q sky130_fd_sc_hd__dfxtp_1
X_15916_ _18407_/CLK _15916_/D vssd1 vssd1 vccd1 vccd1 hold569/A sky130_fd_sc_hd__dfxtp_1
X_11039_ hold2350/X hold5411/X _11153_/C vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16896_ _18067_/CLK _16896_/D vssd1 vssd1 vccd1 vccd1 _16896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ _17715_/CLK _15847_/D vssd1 vssd1 vccd1 vccd1 _15847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _17741_/CLK _15778_/D vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _17517_/CLK _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14729_ hold2409/X _14720_/B _14728_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ _15529_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17448_ _17448_/CLK _17448_/D vssd1 vssd1 vccd1 vccd1 _17448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08181_ _15515_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__or2_1
X_17379_ _17379_/CLK _17379_/D vssd1 vssd1 vccd1 vccd1 _17379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5105 _13687_/X vssd1 vssd1 vccd1 vccd1 _17682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5116 _16548_/Q vssd1 vssd1 vccd1 vccd1 hold5116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5127 _12148_/X vssd1 vssd1 vccd1 vccd1 _17206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_275_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17900_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5138 _16443_/Q vssd1 vssd1 vccd1 vccd1 hold5138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4404 _11314_/X vssd1 vssd1 vccd1 vccd1 _16928_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5149 _10084_/X vssd1 vssd1 vccd1 vccd1 _16518_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4415 hold5824/X vssd1 vssd1 vccd1 vccd1 hold5825/A sky130_fd_sc_hd__buf_4
Xhold4426 _11344_/X vssd1 vssd1 vccd1 vccd1 _16938_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4437 _17635_/Q vssd1 vssd1 vccd1 vccd1 hold4437/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_204_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17891_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4448 _12292_/X vssd1 vssd1 vccd1 vccd1 _17254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3703 _11739_/Y vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4459 _16598_/Q vssd1 vssd1 vccd1 vccd1 hold4459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3714 _11793_/Y vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3725 _16341_/Q vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3736 _10633_/Y vssd1 vssd1 vccd1 vccd1 _16701_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3747 _10624_/Y vssd1 vssd1 vccd1 vccd1 _16698_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3758 _10597_/Y vssd1 vssd1 vccd1 vccd1 _16689_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3769 _12379_/Y vssd1 vssd1 vccd1 vccd1 _17283_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07965_ hold2264/X _07978_/B _07964_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _07965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09704_ hold2263/X _16392_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__mux2_1
X_07896_ _14854_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09635_ hold1389/X hold5425/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__mux2_1
X_09566_ hold1527/X _13238_/A _10271_/S vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08517_ _15521_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _15551_/A _15169_/A hold86/X _15541_/A vssd1 vssd1 vccd1 vccd1 _09498_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_0_182_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08448_ _08504_/A _14913_/A vssd1 vssd1 vccd1 vccd1 _08448_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08379_ _08379_/A hold174/X vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__and2_1
X_10410_ _10524_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ hold1428/X _16954_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__mux2_1
X_10341_ _10551_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ hold4149/X _13059_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
Xhold5650 _11065_/X vssd1 vssd1 vccd1 vccd1 _16845_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10272_ _10491_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__or2_1
Xhold5661 _16835_/Q vssd1 vssd1 vccd1 vccd1 hold5661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5672 _16899_/Q vssd1 vssd1 vccd1 vccd1 hold5672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12011_ hold2014/X _17161_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5683 _16488_/Q vssd1 vssd1 vccd1 vccd1 hold5683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5694 _11572_/X vssd1 vssd1 vccd1 vccd1 _17014_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4960 _13621_/X vssd1 vssd1 vccd1 vccd1 _17660_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4971 _17161_/Q vssd1 vssd1 vccd1 vccd1 hold4971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4982 _12163_/X vssd1 vssd1 vccd1 vccd1 _17211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4993 _17743_/Q vssd1 vssd1 vccd1 vccd1 hold4993/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout460 _13847_/C vssd1 vssd1 vccd1 vccd1 _13859_/C sky130_fd_sc_hd__clkbuf_8
Xfanout471 _11783_/C vssd1 vssd1 vccd1 vccd1 _12329_/C sky130_fd_sc_hd__clkbuf_8
Xfanout482 _11672_/S vssd1 vssd1 vccd1 vccd1 _11219_/C sky130_fd_sc_hd__clkbuf_8
X_16750_ _18337_/CLK _16750_/D vssd1 vssd1 vccd1 vccd1 _16750_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout493 _09893_/S vssd1 vssd1 vccd1 vccd1 _10028_/C sky130_fd_sc_hd__clkbuf_4
X_13962_ hold949/X _13992_/B vssd1 vssd1 vccd1 vccd1 _13962_/X sky130_fd_sc_hd__or2_1
X_15701_ _17777_/CLK _15701_/D vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_79_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17524_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ hold2348/X hold3228/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__mux2_1
X_16681_ _18315_/CLK _16681_/D vssd1 vssd1 vccd1 vccd1 _16681_/Q sky130_fd_sc_hd__dfxtp_1
X_13893_ hold281/A hold242/X vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__nand2_1
X_18420_ _18420_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
X_15632_ _17227_/CLK _15632_/D vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ hold2205/X _17459_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18383_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
X_15563_ _17211_/CLK _15563_/D vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775_ hold2928/X hold3448/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12775_/X sky130_fd_sc_hd__mux2_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/CLK _17302_/D vssd1 vssd1 vccd1 vccd1 _17302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ hold2992/X _14554_/A2 _14513_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14514_/X
+ sky130_fd_sc_hd__o211a_1
X_18282_ _18382_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _17066_/Q _11726_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__and3_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15498_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__and2_1
XFILLER_0_138_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17233_ _17900_/CLK _17233_/D vssd1 vssd1 vccd1 vccd1 _17233_/Q sky130_fd_sc_hd__dfxtp_1
X_14445_ _14786_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14445_/X sky130_fd_sc_hd__or2_1
X_11657_ hold2783/X hold5342/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ hold3678/X _10542_/A _10607_/X vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__a21oi_1
X_17164_ _17260_/CLK _17164_/D vssd1 vssd1 vccd1 vccd1 _17164_/Q sky130_fd_sc_hd__dfxtp_1
X_14376_ _14376_/A hold276/X vssd1 vssd1 vccd1 vccd1 _17987_/D sky130_fd_sc_hd__and2_1
X_11588_ _17868_/Q hold3440/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16115_ _17314_/CLK _16115_/D vssd1 vssd1 vccd1 vccd1 hold528/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold908 hold908/A vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ hold4907/X _13805_/B _13326_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13327_/X
+ sky130_fd_sc_hd__o211a_1
X_17095_ _17221_/CLK _17095_/D vssd1 vssd1 vccd1 vccd1 _17095_/Q sky130_fd_sc_hd__dfxtp_1
Xhold919 hold919/A vssd1 vssd1 vccd1 vccd1 hold919/X sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ _11103_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16096_/CLK _16046_/D vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__dfxtp_1
X_13258_ _17583_/Q _17117_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13258_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ hold2137/X hold3366/X _12308_/C vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__mux2_1
X_13189_ _13188_/X hold3132/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13189_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2309 _14263_/X vssd1 vssd1 vccd1 vccd1 _17932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1608 _15616_/Q vssd1 vssd1 vccd1 vccd1 hold1608/X sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _18061_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1619 _16179_/Q vssd1 vssd1 vccd1 vccd1 hold1619/X sky130_fd_sc_hd__dlygate4sd3_1
X_16948_ _17862_/CLK _16948_/D vssd1 vssd1 vccd1 vccd1 _16948_/Q sky130_fd_sc_hd__dfxtp_1
X_16879_ _18052_/CLK _16879_/D vssd1 vssd1 vccd1 vccd1 _16879_/Q sky130_fd_sc_hd__dfxtp_1
X_09420_ _09438_/B _16296_/Q vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _09400_/A _09351_/B _09360_/B vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_158_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ hold5962/X _08336_/A2 _08301_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _08302_/X
+ sky130_fd_sc_hd__o211a_1
X_09282_ _12813_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _16252_/D sky130_fd_sc_hd__and2_1
XFILLER_0_145_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ hold1022/X _08262_/B _08232_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _15515_/A hold1222/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ hold2326/X _08082_/B _08094_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _08095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4201 _13860_/Y vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4212 _10741_/X vssd1 vssd1 vccd1 vccd1 _16737_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4223 _10144_/X vssd1 vssd1 vccd1 vccd1 _16538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4234 _16817_/Q vssd1 vssd1 vccd1 vccd1 hold4234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3500 _17440_/Q vssd1 vssd1 vccd1 vccd1 hold3500/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4245 _11353_/X vssd1 vssd1 vccd1 vccd1 _16941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4256 _17559_/Q vssd1 vssd1 vccd1 vccd1 hold4256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3511 _17418_/Q vssd1 vssd1 vccd1 vccd1 hold3511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4267 _17254_/Q vssd1 vssd1 vccd1 vccd1 hold4267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3522 _11875_/X vssd1 vssd1 vccd1 vccd1 _17115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3533 _16586_/Q vssd1 vssd1 vccd1 vccd1 hold3533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4278 _11506_/X vssd1 vssd1 vccd1 vccd1 _16992_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3544 _10465_/X vssd1 vssd1 vccd1 vccd1 _16645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4289 _17037_/Q vssd1 vssd1 vccd1 vccd1 hold4289/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2810 _14247_/X vssd1 vssd1 vccd1 vccd1 _17924_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3555 _10372_/X vssd1 vssd1 vccd1 vccd1 _16614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3566 _17703_/Q vssd1 vssd1 vccd1 vccd1 hold3566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 _08235_/X vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 _18143_/Q vssd1 vssd1 vccd1 vccd1 hold2832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3577 _17639_/Q vssd1 vssd1 vccd1 vccd1 hold3577/X sky130_fd_sc_hd__dlygate4sd3_1
X_08997_ hold291/X hold534/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__mux2_1
Xhold2843 _08243_/X vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3588 _17364_/Q vssd1 vssd1 vccd1 vccd1 hold3588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3599 _10002_/Y vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2854 _15730_/Q vssd1 vssd1 vccd1 vccd1 hold2854/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2865 _12671_/X vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2876 _14827_/X vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07948_ _14511_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07948_/X sky130_fd_sc_hd__or2_1
Xhold2887 _17999_/Q vssd1 vssd1 vccd1 vccd1 hold2887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2898 _14747_/X vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07879_ _15557_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__or2_1
X_09618_ _09948_/A _09618_/B vssd1 vssd1 vccd1 vccd1 _09618_/X sky130_fd_sc_hd__or2_1
X_10890_ _11082_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__or2_1
X_09549_ _09933_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ hold3575/X _12559_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _12153_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_197_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18053_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ hold140/X _12509_/A2 _12505_/A3 _12490_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold141/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _14980_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14230_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18355_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11442_ _11637_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ hold871/X _14148_/B _14160_/X _14356_/A vssd1 vssd1 vccd1 vccd1 hold872/A
+ sky130_fd_sc_hd__o211a_1
X_11373_ _11667_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13112_ _13105_/X _13111_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17532_/D sky130_fd_sc_hd__o21a_1
X_10324_ hold4018/X _10646_/B _10323_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10324_/X
+ sky130_fd_sc_hd__o211a_1
X_14092_ _15545_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5480 _16773_/Q vssd1 vssd1 vccd1 vccd1 hold5480/X sky130_fd_sc_hd__dlygate4sd3_1
X_13043_ _13046_/A _13053_/A _13043_/C vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__or3_1
X_10255_ hold4305/X _10619_/B _10254_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _17984_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5491 _10672_/X vssd1 vssd1 vccd1 vccd1 _16714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4790 _15472_/X vssd1 vssd1 vccd1 vccd1 _15473_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17851_ _17884_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_1
X_10186_ hold3487/X _10568_/B _10185_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10186_/X
+ sky130_fd_sc_hd__o211a_1
X_16802_ _18069_/CLK _16802_/D vssd1 vssd1 vccd1 vccd1 _16802_/Q sky130_fd_sc_hd__dfxtp_1
X_17782_ _17877_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
X_14994_ _15209_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__or2_1
Xfanout290 _11115_/A vssd1 vssd1 vccd1 vccd1 _11667_/A sky130_fd_sc_hd__clkbuf_4
X_16733_ _18025_/CLK _16733_/D vssd1 vssd1 vccd1 vccd1 _16733_/Q sky130_fd_sc_hd__dfxtp_1
X_13945_ _15498_/A _13945_/B vssd1 vssd1 vccd1 vccd1 _17780_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16664_ _18222_/CLK _16664_/D vssd1 vssd1 vccd1 vccd1 _16664_/Q sky130_fd_sc_hd__dfxtp_1
X_13876_ _13888_/A _13876_/B vssd1 vssd1 vccd1 vccd1 _13876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18403_ _18410_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
X_15615_ _17211_/CLK _15615_/D vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ hold3054/X _12826_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__mux2_1
X_16595_ _18185_/CLK _16595_/D vssd1 vssd1 vccd1 vccd1 _16595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ _18334_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ hold2062/X _15547_/B _15545_/Y _12885_/A vssd1 vssd1 vccd1 vccd1 _15546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12758_ hold3476/X _12757_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18265_ _18265_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
X_11709_ _12093_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__or2_1
X_15477_ _07805_/A _15477_/A2 _09365_/B hold508/X vssd1 vssd1 vccd1 vccd1 _15480_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12689_ hold3056/X _12688_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17216_ _17216_/CLK _17216_/D vssd1 vssd1 vccd1 vccd1 _17216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ hold2161/X _14433_/B _14427_/Y _14368_/A vssd1 vssd1 vccd1 vccd1 _14428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18196_ _18228_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17147_ _17211_/CLK _17147_/D vssd1 vssd1 vccd1 vccd1 _17147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 hold705/A vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14359_ _14986_/A hold2297/X hold275/X vssd1 vssd1 vccd1 vccd1 _14360_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold716 hold716/A vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold738 la_data_in[20] vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/A vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
X_17078_ _18064_/CLK _17078_/D vssd1 vssd1 vccd1 vccd1 _17078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_13__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_40_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_16029_ _17289_/CLK _16029_/D vssd1 vssd1 vccd1 vccd1 hold446/A sky130_fd_sc_hd__dfxtp_1
X_08920_ hold50/X hold529/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2106 _15599_/Q vssd1 vssd1 vccd1 vccd1 hold2106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2117 _18318_/Q vssd1 vssd1 vccd1 vccd1 hold2117/X sky130_fd_sc_hd__dlygate4sd3_1
X_08851_ _15482_/A _08851_/B vssd1 vssd1 vccd1 vccd1 _16044_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2128 _13981_/X vssd1 vssd1 vccd1 vccd1 _17797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 _18115_/Q vssd1 vssd1 vccd1 vccd1 hold2139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1405 _15660_/Q vssd1 vssd1 vccd1 vccd1 hold1405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _16153_/Q vssd1 vssd1 vccd1 vccd1 hold1416/X sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ _09339_/B _07802_/B vssd1 vssd1 vccd1 vccd1 _07802_/Y sky130_fd_sc_hd__nand2_1
Xhold1427 _08190_/X vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ _15473_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _16011_/D sky130_fd_sc_hd__and2_1
Xhold1438 _18085_/Q vssd1 vssd1 vccd1 vccd1 hold1438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1449 la_data_in[13] vssd1 vssd1 vccd1 vccd1 hold539/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09403_ _07785_/Y hold1504/X _11155_/A vssd1 vssd1 vccd1 vccd1 _16287_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09334_ hold2594/X _09338_/A2 _09333_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09265_ hold265/A _16244_/Q _09277_/S vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_290_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17260_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ hold2091/X _08213_/B _08215_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ _15525_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08078_ _15537_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__or2_1
Xhold4020 _16942_/Q vssd1 vssd1 vccd1 vccd1 hold4020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4031 _10243_/X vssd1 vssd1 vccd1 vccd1 _16571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4042 _13876_/Y vssd1 vssd1 vccd1 vccd1 _17745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4053 _17085_/Q vssd1 vssd1 vccd1 vccd1 hold4053/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4064 _09652_/X vssd1 vssd1 vccd1 vccd1 _16374_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3330 _17466_/Q vssd1 vssd1 vccd1 vccd1 hold3330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4075 _17073_/Q vssd1 vssd1 vccd1 vccd1 hold4075/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3341 _12007_/X vssd1 vssd1 vccd1 vccd1 _17159_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10040_ _16504_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10040_/X sky130_fd_sc_hd__and3_1
Xhold4086 _10549_/X vssd1 vssd1 vccd1 vccd1 _16673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3352 _11617_/X vssd1 vssd1 vccd1 vccd1 _17029_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4097 _16706_/Q vssd1 vssd1 vccd1 vccd1 hold4097/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3363 _11866_/X vssd1 vssd1 vccd1 vccd1 _17112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3374 _11077_/X vssd1 vssd1 vccd1 vccd1 _16849_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__clkbuf_4
Xhold2640 _08222_/X vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3385 _12707_/X vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3396 _17595_/Q vssd1 vssd1 vccd1 vccd1 hold3396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2651 _07897_/X vssd1 vssd1 vccd1 vccd1 _15592_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2662 _16211_/Q vssd1 vssd1 vccd1 vccd1 hold2662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__buf_4
Xhold2673 _15152_/X vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2684 _14593_/X vssd1 vssd1 vccd1 vccd1 _18090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 _16212_/Q vssd1 vssd1 vccd1 vccd1 hold1950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2695 _18457_/Q vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1961 _07872_/X vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _13749_/A _11991_/B vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__or2_1
Xhold1972 _08336_/X vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1983 _15661_/Q vssd1 vssd1 vccd1 vccd1 hold1983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13730_ hold2987/X _17697_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13731_/B sky130_fd_sc_hd__mux2_1
Xhold1994 _16222_/Q vssd1 vssd1 vccd1 vccd1 hold1994/X sky130_fd_sc_hd__dlygate4sd3_1
X_10942_ hold3208/X _11171_/B _10941_/X _14418_/C1 vssd1 vssd1 vccd1 vccd1 _10942_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ hold2772/X _17674_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10873_ hold4488/X _09992_/B _10872_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _10873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15400_ hold548/X _09367_/A _09392_/A hold650/X vssd1 vssd1 vccd1 vccd1 _15400_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ _12927_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _17380_/D sky130_fd_sc_hd__and2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _18315_/CLK _16380_/D vssd1 vssd1 vccd1 vccd1 _16380_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_307_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _15784_/Q hold5110/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _16297_/Q _15477_/A2 _15487_/B1 hold456/X _15330_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12933_/A _12543_/B vssd1 vssd1 vccd1 vccd1 _17357_/D sky130_fd_sc_hd__and2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18050_ _18050_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _15489_/A _15262_/B _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_152_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12474_ _17330_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17001_ _17882_/CLK _17001_/D vssd1 vssd1 vccd1 vccd1 _17001_/Q sky130_fd_sc_hd__dfxtp_1
X_14213_ hold2758/X _14198_/B _14212_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _14213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ hold4555/X _12305_/B _11424_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _15193_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__or2_1
XANTENNA_7 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14144_ _15543_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11356_ hold4087/X _11747_/B _11355_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ hold2744/X hold4675/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__mux2_1
X_14075_ hold1351/X _14105_/A2 _14074_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14075_/X
+ sky130_fd_sc_hd__o211a_1
X_11287_ hold5711/X _11765_/B _11286_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__o211a_1
X_13026_ _17518_/Q hold901/X _13043_/C vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18380_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17903_ _17903_/CLK hold916/X vssd1 vssd1 vccd1 vccd1 hold915/A sky130_fd_sc_hd__dfxtp_1
X_10238_ hold1440/X hold4222/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10239_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18431_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10169_ hold1811/X hold3126/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__mux2_1
X_17834_ _17892_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17765_ _17829_/CLK _17765_/D vssd1 vssd1 vccd1 vccd1 _17765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14977_ hold5959/X _15006_/B hold491/X _15394_/A vssd1 vssd1 vccd1 vccd1 hold492/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13928_ hold235/X _17772_/Q hold244/X vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__mux2_1
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _18241_/CLK _16716_/D vssd1 vssd1 vccd1 vccd1 _16716_/Q sky130_fd_sc_hd__dfxtp_1
X_17696_ _17728_/CLK _17696_/D vssd1 vssd1 vccd1 vccd1 _17696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16647_ _18205_/CLK _16647_/D vssd1 vssd1 vccd1 vccd1 _16647_/Q sky130_fd_sc_hd__dfxtp_1
X_13859_ _17740_/Q _13859_/B _13859_/C vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _18220_/CLK _16578_/D vssd1 vssd1 vccd1 vccd1 _16578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18317_ _18382_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15529_ _15529_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09050_ hold50/X hold247/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__mux2_1
X_18248_ _18416_/CLK hold367/X vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ _14850_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18179_ _18268_/CLK hold767/X vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 hold80/X vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold513/A vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 hold524/A vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold535 hold535/A vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold546 input14/X vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold557 hold557/A vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold568 hold568/A vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09952_ hold5076/X _09952_/A2 _09951_/X _15144_/C1 vssd1 vssd1 vccd1 vccd1 _09952_/X
+ sky130_fd_sc_hd__o211a_1
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08903_ _08970_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _16069_/D sky130_fd_sc_hd__and2_1
X_09883_ hold5140/X _10073_/B _09882_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09883_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _14017_/X vssd1 vssd1 vccd1 vccd1 _17814_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ hold179/X hold307/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__mux2_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _14713_/X vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _15552_/X vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 _17788_/Q vssd1 vssd1 vccd1 vccd1 hold1235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _18357_/Q vssd1 vssd1 vccd1 vccd1 hold1246/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1257 _15680_/Q vssd1 vssd1 vccd1 vccd1 hold1257/X sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ hold184/X hold687/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1268 _15162_/X vssd1 vssd1 vccd1 vccd1 _18364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _08010_/X vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _12438_/A _08696_/B vssd1 vssd1 vccd1 vccd1 _15969_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _15105_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _12777_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _16235_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ hold207/X _15508_/B vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__or2_2
XFILLER_0_105_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _16894_/Q _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11210_/X sky130_fd_sc_hd__and3_1
XFILLER_0_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ hold5001/X _12311_/B _12189_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _12190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11141_ _16871_/Q _11150_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__and3_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput77 _13169_/A vssd1 vssd1 vccd1 vccd1 output77/X sky130_fd_sc_hd__buf_6
X_11072_ hold2866/X hold3194/X _11171_/C vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__mux2_1
Xoutput88 _13249_/A vssd1 vssd1 vccd1 vccd1 output88/X sky130_fd_sc_hd__buf_6
XFILLER_0_179_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput99 _13097_/A vssd1 vssd1 vccd1 vccd1 output99/X sky130_fd_sc_hd__buf_6
Xhold3160 _13824_/Y vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3171 _16353_/Q vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10023_ _13174_/A _09981_/A _10022_/X vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__a21oi_1
X_14900_ _14970_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__or2_1
X_15880_ _17719_/CLK _15880_/D vssd1 vssd1 vccd1 vccd1 _15880_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3182 _16903_/Q vssd1 vssd1 vccd1 vccd1 hold3182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3193 _12355_/Y vssd1 vssd1 vccd1 vccd1 _17275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2470 _08089_/X vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2481 _18439_/Q vssd1 vssd1 vccd1 vccd1 hold2481/X sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ hold960/X _14828_/B _14830_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 hold961/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 _14414_/X vssd1 vssd1 vccd1 vccd1 _18005_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _18185_/CLK _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1780 _18428_/Q vssd1 vssd1 vccd1 vccd1 hold1780/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1791 _14484_/X vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ _15209_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14762_/X sky130_fd_sc_hd__or2_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ hold4599/X _13871_/B _11973_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11974_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _18382_/CLK _16501_/D vssd1 vssd1 vccd1 vccd1 _16501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13713_/A _13713_/B vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _17484_/CLK _17481_/D vssd1 vssd1 vccd1 vccd1 _17481_/Q sky130_fd_sc_hd__dfxtp_1
X_10925_ hold2949/X hold5407/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__mux2_1
X_14693_ hold3029/X _14720_/B _14692_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14693_/X
+ sky130_fd_sc_hd__o211a_1
X_16432_ _18391_/CLK _16432_/D vssd1 vssd1 vccd1 vccd1 _16432_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_141_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13644_ _13776_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10856_ hold2297/X hold4371/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _18308_/CLK _16363_/D vssd1 vssd1 vccd1 vccd1 _16363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13767_/A _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__or2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ hold1443/X _16753_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10788_/B sky130_fd_sc_hd__mux2_1
X_18102_ _18232_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__and2_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ hold1420/X _17353_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__mux2_1
X_16294_ _16314_/CLK _16294_/D vssd1 vssd1 vccd1 vccd1 _16294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18033_ _18033_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
X_15245_ hold424/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__or2_1
X_12457_ hold41/X _12509_/A2 _12505_/A3 _12456_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold42/A sky130_fd_sc_hd__o311a_1
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ hold1035/X _16960_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__mux2_1
X_15176_ hold958/X hold609/X _15175_/X _15394_/A vssd1 vssd1 vccd1 vccd1 hold959/A
+ sky130_fd_sc_hd__o211a_1
X_12388_ _15374_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _17287_/D sky130_fd_sc_hd__and2_1
X_14127_ hold2609/X _14148_/B _14126_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__o211a_1
X_11339_ hold1561/X hold4455/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ hold756/X _14072_/B vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _14972_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__or2_1
X_17817_ _17884_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_1
X_08550_ hold443/X hold558/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08551_/B sky130_fd_sc_hd__mux2_1
X_17748_ _17748_/CLK _17748_/D vssd1 vssd1 vccd1 vccd1 _17748_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_229_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17282_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08481_ hold1445/X _08486_/B _08480_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08481_/X
+ sky130_fd_sc_hd__o211a_1
X_17679_ _17743_/CLK _17679_/D vssd1 vssd1 vccd1 vccd1 _17679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ _15543_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _15414_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _16133_/D sky130_fd_sc_hd__and2_1
XFILLER_0_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold332 la_data_in[18] vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold343 input10/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold489/X vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__buf_6
Xhold376 hold376/A vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 hold387/A vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout801 _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14831_/C1 sky130_fd_sc_hd__buf_4
X_09935_ hold1290/X hold5371/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__mux2_1
Xfanout812 fanout816/X vssd1 vssd1 vccd1 vccd1 _15144_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout823 _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__buf_4
Xfanout834 fanout841/X vssd1 vssd1 vccd1 vccd1 _14955_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout845 _11791_/A vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__clkbuf_8
Xfanout856 _17754_/Q vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__buf_12
Xfanout867 _07782_/Y vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__buf_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ hold2672/X hold4329/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__mux2_1
Xhold1010 _15829_/Q vssd1 vssd1 vccd1 vccd1 hold1010/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 _15199_/A vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__clkbuf_16
Xhold1021 _14577_/X vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 _14854_/A vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__buf_6
XFILLER_0_175_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08817_ _15491_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _16027_/D sky130_fd_sc_hd__and2_1
Xhold1032 _08388_/X vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _17889_/Q vssd1 vssd1 vccd1 vccd1 hold1043/X sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ hold2159/X _16423_/Q _09893_/S vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__mux2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _14411_/X vssd1 vssd1 vccd1 vccd1 hold1054/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _17796_/Q vssd1 vssd1 vccd1 vccd1 hold1065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 _09069_/X vssd1 vssd1 vccd1 vccd1 _16149_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _15414_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _15994_/D sky130_fd_sc_hd__and2_1
Xhold1087 _15809_/Q vssd1 vssd1 vccd1 vccd1 hold1087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 hold1098/A vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__buf_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ hold47/X hold580/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__mux2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _11121_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ hold2230/X hold4099/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ hold3728/X _10554_/A _10640_/X vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ hold4783/X _13868_/B _13359_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13360_/X
+ sky130_fd_sc_hd__o211a_1
X_10572_ hold3662/X _10380_/A _10571_/X vssd1 vssd1 vccd1 vccd1 _10572_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ _17261_/Q _12311_/B _13793_/S vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13291_ _13290_/X hold5902/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15030_ _15030_/A _15030_/B vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ hold2220/X _17238_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ hold2106/X hold4482/X _13844_/C vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _11670_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or2_1
X_16981_ _17829_/CLK _16981_/D vssd1 vssd1 vccd1 vccd1 _16981_/Q sky130_fd_sc_hd__dfxtp_1
X_15932_ _17530_/CLK _15932_/D vssd1 vssd1 vccd1 vccd1 hold601/A sky130_fd_sc_hd__dfxtp_1
X_11055_ _11061_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__or2_1
X_10006_ _11203_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10006_/Y sky130_fd_sc_hd__nor2_1
X_15863_ _17736_/CLK _15863_/D vssd1 vssd1 vccd1 vccd1 _15863_/Q sky130_fd_sc_hd__dfxtp_1
X_14814_ _15099_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17602_ _17634_/CLK _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
X_15794_ _17725_/CLK _15794_/D vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_322_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17754_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _18308_/CLK _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_1
X_14745_ hold1344/X _14772_/B _14744_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14745_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11957_ hold837/X hold4795/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17464_ _17464_/CLK _17464_/D vssd1 vssd1 vccd1 vccd1 _17464_/Q sky130_fd_sc_hd__dfxtp_1
X_10908_ _11097_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__or2_1
X_14676_ _15231_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14676_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11888_ hold1308/X hold3147/X _12368_/C vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16415_ _18392_/CLK _16415_/D vssd1 vssd1 vccd1 vccd1 _16415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13627_ hold4500/X _13814_/B _13626_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _13627_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17395_ _18448_/CLK _17395_/D vssd1 vssd1 vccd1 vccd1 _17395_/Q sky130_fd_sc_hd__dfxtp_1
X_10839_ _11031_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16346_ _18355_/CLK _16346_/D vssd1 vssd1 vccd1 vccd1 _16346_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ hold3579/X _13886_/B _13557_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12509_ hold38/X _12509_/A2 _12445_/B _12508_/X _09021_/A vssd1 vssd1 vccd1 vccd1
+ hold39/A sky130_fd_sc_hd__o311a_1
XFILLER_0_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16277_ _17379_/CLK _16277_/D vssd1 vssd1 vccd1 vccd1 _16277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ hold4816/X _13868_/B _13488_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13489_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5309 _16731_/Q vssd1 vssd1 vccd1 vccd1 hold5309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ hold2756/X _15219_/B _15227_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15228_/X
+ sky130_fd_sc_hd__o211a_1
X_18016_ _18305_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4608 _09751_/X vssd1 vssd1 vccd1 vccd1 _16407_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4619 _16936_/Q vssd1 vssd1 vccd1 vccd1 hold4619/X sky130_fd_sc_hd__dlygate4sd3_1
X_15159_ _15213_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__or2_1
Xhold3907 _17561_/Q vssd1 vssd1 vccd1 vccd1 hold3907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3918 _09625_/X vssd1 vssd1 vccd1 vccd1 _16365_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3929 _16873_/Q vssd1 vssd1 vccd1 vccd1 hold3929/X sky130_fd_sc_hd__dlygate4sd3_1
X_07981_ hold1826/X _07978_/B _07980_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _07981_/X
+ sky130_fd_sc_hd__o211a_1
X_09720_ _09924_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__or2_1
X_09651_ _10380_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ _15374_/A _08602_/B vssd1 vssd1 vccd1 vccd1 _15923_/D sky130_fd_sc_hd__and2_1
X_09582_ _10098_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08533_ _15244_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _15890_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08464_ _14517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _14218_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5810 hold5931/X vssd1 vssd1 vccd1 vccd1 _13137_/A sky130_fd_sc_hd__dlygate4sd3_1
X_09016_ hold126/X hold700/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5821 hold5821/A vssd1 vssd1 vccd1 vccd1 load_status[0] sky130_fd_sc_hd__buf_12
Xhold5832 _17523_/Q vssd1 vssd1 vccd1 vccd1 hold5832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5843 hold5843/A vssd1 vssd1 vccd1 vccd1 hold5843/X sky130_fd_sc_hd__buf_2
Xhold5854 hold5941/X vssd1 vssd1 vccd1 vccd1 hold5854/X sky130_fd_sc_hd__clkbuf_2
Xhold140 hold480/X vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__clkbuf_4
Xhold5865 hold5865/A vssd1 vssd1 vccd1 vccd1 hold5865/X sky130_fd_sc_hd__buf_2
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5876 hold5983/X vssd1 vssd1 vccd1 vccd1 hold5876/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold162 input6/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__clkbuf_8
Xhold5887 _09483_/X vssd1 vssd1 vccd1 vccd1 hold5887/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold5898 _16920_/Q vssd1 vssd1 vccd1 vccd1 hold5898/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold412/X vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__buf_4
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__buf_1
Xfanout620 _15486_/A2 vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkbuf_8
Xfanout631 _07824_/Y vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__clkbuf_4
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__or2_1
Xfanout642 _12810_/A vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__buf_4
Xfanout653 fanout660/X vssd1 vssd1 vccd1 vccd1 _12927_/A sky130_fd_sc_hd__buf_2
Xfanout664 fanout842/X vssd1 vssd1 vccd1 vccd1 _13627_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14149_/C1 sky130_fd_sc_hd__buf_4
Xfanout686 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__buf_2
Xfanout697 _08585_/A vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__clkbuf_4
X_09849_ _11082_/A _09849_/B vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__or2_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ hold3309/X _12859_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__mux2_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11811_ _13797_/A _11811_/B vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ hold3500/X _12790_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ hold1727/X _14541_/B _14529_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14530_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ hold3156/X _11649_/A _11741_/X vssd1 vssd1 vccd1 vccd1 _11742_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ _14980_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14461_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11697_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__or2_1
XFILLER_0_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16200_ _17484_/CLK _16200_/D vssd1 vssd1 vccd1 vccd1 _16200_/Q sky130_fd_sc_hd__dfxtp_1
X_13412_ hold2431/X hold3313/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10624_ _10651_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10624_/Y sky130_fd_sc_hd__nor2_1
X_17180_ _17584_/CLK _17180_/D vssd1 vssd1 vccd1 vccd1 _17180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14392_ _14392_/A _14392_/B vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__and2_1
X_16131_ _18413_/CLK _16131_/D vssd1 vssd1 vccd1 vccd1 hold670/A sky130_fd_sc_hd__dfxtp_1
X_13343_ hold1644/X hold3159/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10555_ hold4065/X _10640_/B _10554_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _17513_/CLK _16062_/D vssd1 vssd1 vccd1 vccd1 hold564/A sky130_fd_sc_hd__dfxtp_1
X_13274_ _17585_/Q _17119_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ hold4287/X _10580_/B _10485_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ hold2532/X _15004_/B _15012_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _13794_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__or2_1
X_12156_ _12255_/A _12156_/B vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__or2_1
X_11107_ hold5627/X _11201_/B _11106_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _11107_/X
+ sky130_fd_sc_hd__o211a_1
X_12087_ _13749_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16964_ _18427_/CLK _16964_/D vssd1 vssd1 vccd1 vccd1 _16964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15915_ _17313_/CLK _15915_/D vssd1 vssd1 vccd1 vccd1 hold522/A sky130_fd_sc_hd__dfxtp_1
X_11038_ hold5558/X _09992_/B _11037_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _11038_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _18190_/CLK _16895_/D vssd1 vssd1 vccd1 vccd1 _16895_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _17649_/CLK hold846/X vssd1 vssd1 vccd1 vccd1 hold845/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _17740_/CLK _15777_/D vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfxtp_1
X_12989_ hold3418/X _12988_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__mux2_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17516_ _17516_/CLK _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14728_ _14728_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__or2_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ hold1191/X _14664_/B _14658_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14659_/X
+ sky130_fd_sc_hd__o211a_1
X_17447_ _17447_/CLK _17447_/D vssd1 vssd1 vccd1 vccd1 _17447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08180_ hold2987/X _08209_/B _08179_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08180_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17378_ _17379_/CLK _17378_/D vssd1 vssd1 vccd1 vccd1 _17378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16329_ _18243_/CLK _16329_/D vssd1 vssd1 vccd1 vccd1 _16329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5106 _17149_/Q vssd1 vssd1 vccd1 vccd1 hold5106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5117 _10078_/X vssd1 vssd1 vccd1 vccd1 _16516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5128 _17135_/Q vssd1 vssd1 vccd1 vccd1 hold5128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5139 _09763_/X vssd1 vssd1 vccd1 vccd1 _16411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4405 _16829_/Q vssd1 vssd1 vccd1 vccd1 hold4405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4416 _15343_/X vssd1 vssd1 vccd1 vccd1 _15344_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4427 _17093_/Q vssd1 vssd1 vccd1 vccd1 hold4427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4438 _13450_/X vssd1 vssd1 vccd1 vccd1 _17603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4449 _16668_/Q vssd1 vssd1 vccd1 vccd1 hold4449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3704 _11740_/Y vssd1 vssd1 vccd1 vccd1 _17070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3715 _11794_/Y vssd1 vssd1 vccd1 vccd1 _17088_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3726 _10032_/Y vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3737 _16907_/Q vssd1 vssd1 vccd1 vccd1 hold3737/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3748 hold4479/X vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3759 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold3759/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_244_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17740_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07964_ _15533_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09703_ hold5612/X _10022_/B _09702_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _09703_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07895_ hold1142/X _07918_/B _07894_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07895_/X
+ sky130_fd_sc_hd__o211a_1
X_09634_ hold5635/X _11201_/B _09633_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _09634_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09565_ hold3386/X _10049_/B _09564_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ hold1838/X _08503_/Y _08515_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _08516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09496_ _09496_/A hold799/X hold770/X vssd1 vssd1 vccd1 vccd1 _09498_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ hold279/X hold298/A hold606/A hold624/A vssd1 vssd1 vccd1 vccd1 _14913_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_93_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08378_ hold173/X _15821_/Q hold122/X vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__mux2_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10340_ hold2846/X hold3326/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5640 _09544_/X vssd1 vssd1 vccd1 vccd1 _16338_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10271_ hold2959/X _16581_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__mux2_1
Xhold5651 _16897_/Q vssd1 vssd1 vccd1 vccd1 hold5651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5662 _16866_/Q vssd1 vssd1 vccd1 vccd1 hold5662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5673 _11131_/X vssd1 vssd1 vccd1 vccd1 _16867_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12010_ hold4739/X _13811_/B _12009_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _12010_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5684 _09898_/X vssd1 vssd1 vccd1 vccd1 _16456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4950 _13792_/X vssd1 vssd1 vccd1 vccd1 _17717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5695 _16388_/Q vssd1 vssd1 vccd1 vccd1 hold5695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4961 _17276_/Q vssd1 vssd1 vccd1 vccd1 hold4961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4972 _11917_/X vssd1 vssd1 vccd1 vccd1 _17129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4983 _17732_/Q vssd1 vssd1 vccd1 vccd1 hold4983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4994 _13774_/X vssd1 vssd1 vccd1 vccd1 _17711_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout450 _11717_/C vssd1 vssd1 vccd1 vccd1 _11726_/C sky130_fd_sc_hd__clkbuf_8
Xfanout461 fanout484/X vssd1 vssd1 vccd1 vccd1 _13847_/C sky130_fd_sc_hd__buf_4
Xfanout472 _11783_/C vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__clkbuf_8
X_13961_ hold2769/X _13980_/B _13960_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _13961_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout483 fanout484/X vssd1 vssd1 vccd1 vccd1 _11672_/S sky130_fd_sc_hd__buf_4
Xfanout494 _10763_/S vssd1 vssd1 vccd1 vccd1 _09893_/S sky130_fd_sc_hd__clkbuf_4
X_15700_ _17268_/CLK _15700_/D vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfxtp_1
X_12912_ _12918_/A _12912_/B vssd1 vssd1 vccd1 vccd1 _17480_/D sky130_fd_sc_hd__and2_1
X_16680_ _18205_/CLK _16680_/D vssd1 vssd1 vccd1 vccd1 _16680_/Q sky130_fd_sc_hd__dfxtp_1
X_13892_ hold241/X hold271/X vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__or2_1
X_12843_ _12843_/A _12843_/B vssd1 vssd1 vccd1 vccd1 _17457_/D sky130_fd_sc_hd__and2_1
X_15631_ _17227_/CLK _15631_/D vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _18381_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15562_ _17275_/CLK _15562_/D vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12777_/A _12774_/B vssd1 vssd1 vccd1 vccd1 _17434_/D sky130_fd_sc_hd__and2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17307_/CLK _17301_/D vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _15193_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _12301_/A _11725_/B vssd1 vssd1 vccd1 vccd1 _11725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15493_ _14218_/A hold1767/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15494_/B sky130_fd_sc_hd__mux2_1
X_18281_ _18391_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17232_ _17232_/CLK _17232_/D vssd1 vssd1 vccd1 vccd1 _17232_/Q sky130_fd_sc_hd__dfxtp_1
X_14444_ hold2921/X _14433_/B _14443_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11656_ hold5653/X _12329_/B _11655_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _16693_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__and3_1
X_17163_ _18428_/CLK _17163_/D vssd1 vssd1 vccd1 vccd1 _17163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14375_ hold235/X _17987_/Q hold275/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ hold4538/X _12320_/B _11586_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _17329_/CLK _16114_/D vssd1 vssd1 vccd1 vccd1 hold453/A sky130_fd_sc_hd__dfxtp_1
X_13326_ _13710_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17094_ _17592_/CLK _17094_/D vssd1 vssd1 vccd1 vccd1 _17094_/Q sky130_fd_sc_hd__dfxtp_1
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ hold855/X _16670_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _17307_/CLK _16045_/D vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13257_ _13257_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__and2_1
Xclkbuf_5_12__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_47_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10469_ hold960/X hold4901/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ hold4433/X _13811_/B _12207_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188_ hold3849/X _13187_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12139_ hold5472/X _12329_/B _12138_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _12139_/X
+ sky130_fd_sc_hd__o211a_1
X_17996_ _18208_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1609 _07947_/X vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _17827_/CLK _16947_/D vssd1 vssd1 vccd1 vccd1 _16947_/Q sky130_fd_sc_hd__dfxtp_1
X_16878_ _18062_/CLK _16878_/D vssd1 vssd1 vccd1 vccd1 _16878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15829_ _17725_/CLK _15829_/D vssd1 vssd1 vccd1 vccd1 _15829_/Q sky130_fd_sc_hd__dfxtp_1
X_09350_ _15543_/A _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09360_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_176_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ _15199_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08301_/X sky130_fd_sc_hd__or2_1
X_09281_ _15557_/A hold2710/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08232_ hold756/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08163_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _15719_/D sky130_fd_sc_hd__and2_1
XFILLER_0_172_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08094_ _15553_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4202 _13861_/Y vssd1 vssd1 vccd1 vccd1 _17740_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4213 _16656_/Q vssd1 vssd1 vccd1 vccd1 hold4213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4224 _16578_/Q vssd1 vssd1 vccd1 vccd1 hold4224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4235 _10885_/X vssd1 vssd1 vccd1 vccd1 _16785_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3501 _12791_/X vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4246 _16562_/Q vssd1 vssd1 vccd1 vccd1 hold4246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3512 _17417_/Q vssd1 vssd1 vccd1 vccd1 hold3512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4257 _16804_/Q vssd1 vssd1 vccd1 vccd1 hold4257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4268 _12196_/X vssd1 vssd1 vccd1 vccd1 _17222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3523 _17444_/Q vssd1 vssd1 vccd1 vccd1 hold3523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4279 _16409_/Q vssd1 vssd1 vccd1 vccd1 hold4279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3534 _10192_/X vssd1 vssd1 vccd1 vccd1 _16554_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2800 _14785_/X vssd1 vssd1 vccd1 vccd1 _18183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3545 hold6011/X vssd1 vssd1 vccd1 vccd1 hold3545/X sky130_fd_sc_hd__buf_2
Xhold2811 _15782_/Q vssd1 vssd1 vccd1 vccd1 hold2811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3556 _17679_/Q vssd1 vssd1 vccd1 vccd1 hold3556/X sky130_fd_sc_hd__dlygate4sd3_1
X_08996_ _12442_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _16115_/D sky130_fd_sc_hd__and2_1
Xhold3567 _13654_/X vssd1 vssd1 vccd1 vccd1 _17671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2822 _18008_/Q vssd1 vssd1 vccd1 vccd1 hold2822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 _14703_/X vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3578 _13462_/X vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3589 _12563_/X vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2844 _17929_/Q vssd1 vssd1 vccd1 vccd1 hold2844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 _08188_/X vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07947_ hold1608/X _07991_/A2 _07946_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07947_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2866 _18051_/Q vssd1 vssd1 vccd1 vccd1 hold2866/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2877 _17766_/Q vssd1 vssd1 vccd1 vccd1 hold2877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2888 _14402_/X vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2899 _17927_/Q vssd1 vssd1 vccd1 vccd1 hold2899/X sky130_fd_sc_hd__dlygate4sd3_1
X_07878_ hold2318/X _07865_/B _07877_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _07878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09617_ hold2838/X hold3831/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ hold1220/X _13190_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09479_ hold634/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09481_/C sky130_fd_sc_hd__or2_1
XFILLER_0_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11510_ hold1351/X hold4153/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__mux2_1
X_12490_ _17338_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11441_ hold2616/X hold4611/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ hold784/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__or2_1
X_11372_ hold1065/X _16948_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11373_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _13183_/A1 _13109_/X _13110_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13111_/X
+ sky130_fd_sc_hd__o211a_1
X_10323_ _10521_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14091_ hold1881/X _14094_/B _14090_/Y _15504_/A vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_166_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18206_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13042_ _13046_/C _13046_/D hold794/X vssd1 vssd1 vccd1 vccd1 hold795/A sky130_fd_sc_hd__nor3_1
Xhold5470 _17076_/Q vssd1 vssd1 vccd1 vccd1 hold5470/X sky130_fd_sc_hd__dlygate4sd3_1
X_10254_ _10524_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__or2_1
Xhold5481 _10753_/X vssd1 vssd1 vccd1 vccd1 _16741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5492 _16444_/Q vssd1 vssd1 vccd1 vccd1 hold5492/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4780 _10273_/X vssd1 vssd1 vccd1 vccd1 _16581_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17850_ _17884_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
X_10185_ _10560_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__or2_1
Xhold4791 _16790_/Q vssd1 vssd1 vccd1 vccd1 hold4791/X sky130_fd_sc_hd__dlygate4sd3_1
X_16801_ _18070_/CLK _16801_/D vssd1 vssd1 vccd1 vccd1 _16801_/Q sky130_fd_sc_hd__dfxtp_1
X_17781_ _17877_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_1
X_14993_ hold1389/X _15006_/B _14992_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _14993_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout280 _13779_/A vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__buf_4
Xfanout291 fanout298/X vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16732_ _18060_/CLK _16732_/D vssd1 vssd1 vccd1 vccd1 _16732_/Q sky130_fd_sc_hd__dfxtp_1
X_13944_ _15559_/A hold1947/X hold244/X vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__mux2_1
X_16663_ _18221_/CLK _16663_/D vssd1 vssd1 vccd1 vccd1 _16663_/Q sky130_fd_sc_hd__dfxtp_1
X_13875_ hold4041/X _13791_/A _13874_/X vssd1 vssd1 vccd1 vccd1 _13876_/B sky130_fd_sc_hd__a21oi_1
X_18402_ _18409_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12826_ hold1879/X hold3044/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12826_/X sky130_fd_sc_hd__mux2_1
X_15614_ _17274_/CLK _15614_/D vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _18216_/CLK _16594_/D vssd1 vssd1 vccd1 vccd1 _16594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18333_ _18399_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ hold2290/X hold3122/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__mux2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15545_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ hold2631/X hold4627/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__mux2_1
X_18264_ _18392_/CLK hold862/X vssd1 vssd1 vccd1 vccd1 hold861/A sky130_fd_sc_hd__dfxtp_1
X_15476_ hold257/X _09392_/B _09386_/D hold181/X _15475_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12688_ hold2244/X hold3050/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17215_ _17282_/CLK _17215_/D vssd1 vssd1 vccd1 vccd1 _17215_/Q sky130_fd_sc_hd__dfxtp_1
X_14427_ _15541_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__nand2_1
X_11639_ hold2732/X hold4289/X _11735_/C vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__mux2_1
X_18195_ _18227_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ _17274_/CLK _17146_/D vssd1 vssd1 vccd1 vccd1 _17146_/Q sky130_fd_sc_hd__dfxtp_1
X_14358_ _14360_/A _14358_/B vssd1 vssd1 vccd1 vccd1 _17978_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold706 hold706/A vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _13308_/X hold3126/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold728 hold738/X vssd1 vssd1 vccd1 vccd1 hold739/A sky130_fd_sc_hd__dlygate4sd3_1
X_17077_ _17799_/CLK _17077_/D vssd1 vssd1 vccd1 vccd1 _17077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold739 hold739/A vssd1 vssd1 vccd1 vccd1 input49/A sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ hold1197/X _14333_/A2 _14288_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14289_/X
+ sky130_fd_sc_hd__o211a_1
X_16028_ _17284_/CLK _16028_/D vssd1 vssd1 vccd1 vccd1 hold376/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08850_ hold149/X hold167/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08851_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2107 _07911_/X vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2118 _18266_/Q vssd1 vssd1 vccd1 vccd1 hold2118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2129 _15579_/Q vssd1 vssd1 vccd1 vccd1 hold2129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1406 _08038_/X vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07801_ _09342_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__and2_1
X_08781_ hold50/X hold261/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__mux2_1
Xhold1417 _09077_/X vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 _17802_/Q vssd1 vssd1 vccd1 vccd1 hold1428/X sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _18431_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1439 _14583_/X vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09402_ _15354_/A _09402_/B vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__and2_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09333_ hold800/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _12753_/A hold918/X vssd1 vssd1 vccd1 vccd1 _16243_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _15549_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08215_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ hold1361/X _09216_/B _09194_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _09195_/X
+ sky130_fd_sc_hd__o211a_1
X_08146_ _14330_/A hold1308/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__mux2_1
X_08077_ hold1740/X _08088_/B _08076_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _08077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4010 _16784_/Q vssd1 vssd1 vccd1 vccd1 hold4010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4021 _11260_/X vssd1 vssd1 vccd1 vccd1 _16910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4032 _17560_/Q vssd1 vssd1 vccd1 vccd1 hold4032/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4043 _16876_/Q vssd1 vssd1 vccd1 vccd1 hold4043/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4054 _11689_/X vssd1 vssd1 vccd1 vccd1 _17053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3320 _17130_/Q vssd1 vssd1 vccd1 vccd1 hold3320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4065 _16707_/Q vssd1 vssd1 vccd1 vccd1 hold4065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4076 _11653_/X vssd1 vssd1 vccd1 vccd1 _17041_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3331 _17464_/Q vssd1 vssd1 vccd1 vccd1 hold3331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3342 _16601_/Q vssd1 vssd1 vccd1 vccd1 hold3342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4087 _16974_/Q vssd1 vssd1 vccd1 vccd1 hold4087/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4098 _10552_/X vssd1 vssd1 vccd1 vccd1 _16674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3353 _17166_/Q vssd1 vssd1 vccd1 vccd1 hold3353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3364 _16697_/Q vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkbuf_2
Xhold2630 _15700_/Q vssd1 vssd1 vccd1 vccd1 hold2630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3375 _17375_/Q vssd1 vssd1 vccd1 vccd1 hold3375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3386 _16377_/Q vssd1 vssd1 vccd1 vccd1 hold3386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2641 _18066_/Q vssd1 vssd1 vccd1 vccd1 hold2641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold96/X vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_4
X_08979_ hold140/X hold691/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__mux2_1
Xhold3397 _13330_/X vssd1 vssd1 vccd1 vccd1 _17563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2652 _16225_/Q vssd1 vssd1 vccd1 vccd1 hold2652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2663 _09199_/X vssd1 vssd1 vccd1 vccd1 _16211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2674 _15593_/Q vssd1 vssd1 vccd1 vccd1 hold2674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 _18133_/Q vssd1 vssd1 vccd1 vccd1 hold2685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 _14035_/X vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 _09201_/X vssd1 vssd1 vccd1 vccd1 _16212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ hold1654/X hold4389/X _13844_/C vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__mux2_1
Xhold2696 _15558_/X vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1962 _18367_/Q vssd1 vssd1 vccd1 vccd1 hold1962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1973 _18123_/Q vssd1 vssd1 vccd1 vccd1 hold1973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 _08040_/X vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1995 _09221_/X vssd1 vssd1 vccd1 vccd1 _16222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _11076_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ hold5144/X _13883_/B _13659_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13660_/X
+ sky130_fd_sc_hd__o211a_1
X_10872_ _11067_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__or2_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ hold3346/X _12610_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ hold5092/X _13880_/B _13590_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13591_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ hold553/X _15486_/A2 _15446_/B1 hold564/X vssd1 vssd1 vccd1 vccd1 _15330_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ hold3581/X _12541_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _16290_/Q _15477_/A2 _15487_/B1 hold529/X _15260_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/D sky130_fd_sc_hd__a221o_1
X_12473_ hold59/X _08598_/B _08999_/B _12472_/X _15344_/A vssd1 vssd1 vccd1 vccd1
+ hold60/A sky130_fd_sc_hd__o311a_1
X_17000_ _17880_/CLK _17000_/D vssd1 vssd1 vccd1 vccd1 _17000_/Q sky130_fd_sc_hd__dfxtp_1
X_14212_ _15557_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ _12018_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__or2_1
X_15192_ hold1525/X _15219_/B _15191_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15192_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_8 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14143_ hold2172/X hold587/X _14142_/Y _13943_/A vssd1 vssd1 vccd1 vccd1 _14143_/X
+ sky130_fd_sc_hd__o211a_1
X_11355_ _11652_/A _11355_/B vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10306_ hold4799/X _10646_/B _10305_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10306_/X
+ sky130_fd_sc_hd__o211a_1
X_14074_ hold883/X _14106_/B vssd1 vssd1 vccd1 vccd1 _14074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11286_ _11670_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__or2_1
X_13025_ _13039_/A _13025_/B hold902/X vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__and3_1
X_17902_ _17902_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_1
X_10237_ hold3342/X _10619_/B _10236_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10237_/X
+ sky130_fd_sc_hd__o211a_1
X_17833_ _17892_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_1
X_10168_ hold4224/X _10646_/B _10167_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10168_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _17862_/CLK hold885/X vssd1 vssd1 vccd1 vccd1 _17764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10099_ hold3524/X _10073_/B _10098_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10099_/X
+ sky130_fd_sc_hd__o211a_1
X_14976_ hold490/X _15018_/B vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16715_ _18305_/CLK _16715_/D vssd1 vssd1 vccd1 vccd1 _16715_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_63_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _16314_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13927_ _13929_/A hold245/X vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__and2_1
XFILLER_0_156_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17695_ _17730_/CLK _17695_/D vssd1 vssd1 vccd1 vccd1 _17695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16646_ _18236_/CLK _16646_/D vssd1 vssd1 vccd1 vccd1 _16646_/Q sky130_fd_sc_hd__dfxtp_1
X_13858_ _13873_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_187_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12809_ hold3517/X _12808_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16577_ _18231_/CLK _16577_/D vssd1 vssd1 vccd1 vccd1 _16577_/Q sky130_fd_sc_hd__dfxtp_1
X_13789_ hold5209/X _13883_/B _13788_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _18380_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ hold2548/X _15547_/B _15527_/X _12885_/A vssd1 vssd1 vccd1 vccd1 _15528_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _18424_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ hold451/X _09386_/A _15479_/A2 _17321_/Q _15458_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ hold2860/X _08033_/B _07999_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _08000_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18178_ _18210_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold503 input8/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17129_ _17878_/CLK _17129_/D vssd1 vssd1 vccd1 vccd1 _17129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold525 hold525/A vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold536 hold536/A vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 hold547/A vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 hold558/A vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _09951_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__or2_1
Xhold569 hold569/A vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ hold214/X hold650/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__mux2_1
X_09882_ _10506_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__or2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08833_ _15314_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _16035_/D sky130_fd_sc_hd__and2_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _15702_/Q vssd1 vssd1 vccd1 vccd1 hold1203/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _15617_/Q vssd1 vssd1 vccd1 vccd1 hold1214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 _15862_/Q vssd1 vssd1 vccd1 vccd1 hold1225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1236 _13963_/X vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _15148_/X vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _15334_/A hold215/X vssd1 vssd1 vccd1 vccd1 _16002_/D sky130_fd_sc_hd__and2_1
Xhold1258 _08081_/X vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _15576_/Q vssd1 vssd1 vccd1 vccd1 hold1269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ hold179/X hold239/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08696_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09316_ hold2483/X _09325_/B _09315_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ hold949/X hold1107/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ hold207/X _15508_/B vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ _13939_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _15703_/D sky130_fd_sc_hd__and2_1
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ hold4987/X _11732_/B _11139_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11140_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput78 _13177_/A vssd1 vssd1 vccd1 vccd1 output78/X sky130_fd_sc_hd__buf_6
X_11071_ hold5723/X _11747_/B _11070_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11071_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput89 _13257_/A vssd1 vssd1 vccd1 vccd1 output89/X sky130_fd_sc_hd__buf_6
Xhold3150 _17563_/Q vssd1 vssd1 vccd1 vccd1 hold3150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10022_ _16498_/Q _10022_/B _10022_/C vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__and3_1
Xhold3161 _13825_/Y vssd1 vssd1 vccd1 vccd1 _17728_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3172 _10068_/Y vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3183 _11718_/Y vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3194 _16848_/Q vssd1 vssd1 vccd1 vccd1 hold3194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2460 _15180_/X vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2471 _15647_/Q vssd1 vssd1 vccd1 vccd1 hold2471/X sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ hold730/X _14840_/B vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__or2_1
Xhold2482 _15522_/X vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 _17839_/Q vssd1 vssd1 vccd1 vccd1 hold2493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 hold6002/X vssd1 vssd1 vccd1 vccd1 input1/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14761_ hold2901/X _14772_/B _14760_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _14761_/X
+ sky130_fd_sc_hd__o211a_1
X_11973_ _13392_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__or2_1
Xhold1781 _16267_/Q vssd1 vssd1 vccd1 vccd1 hold1781/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 _15606_/Q vssd1 vssd1 vccd1 vccd1 hold1792/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _18363_/CLK _16500_/D vssd1 vssd1 vccd1 vccd1 _16500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ hold2352/X _17691_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13713_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ hold5484/X _11762_/B _10923_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _10924_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17480_/CLK _17480_/D vssd1 vssd1 vccd1 vccd1 _17480_/Q sky130_fd_sc_hd__dfxtp_1
X_14692_ _15193_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__or2_1
X_16431_ _18381_/CLK _16431_/D vssd1 vssd1 vccd1 vccd1 _16431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13643_ hold1971/X _17668_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__mux2_1
X_10855_ hold4373/X _11726_/B _10854_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _10855_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ hold2997/X _17645_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13575_/B sky130_fd_sc_hd__mux2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _18371_/CLK _16362_/D vssd1 vssd1 vccd1 vccd1 _16362_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ hold4010/X _11747_/B _10785_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _10786_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18223_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15490_/A1 _15305_/X _15312_/X _15490_/B1 hold4867/X vssd1 vssd1 vccd1 vccd1
+ _15313_/X sky130_fd_sc_hd__a32o_1
X_12525_ _13002_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _17351_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _17511_/CLK _16293_/D vssd1 vssd1 vccd1 vccd1 _16293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_181_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18059_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18032_ _18032_/CLK hold821/X vssd1 vssd1 vccd1 vccd1 hold820/A sky130_fd_sc_hd__dfxtp_1
X_12456_ _17321_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__or2_1
X_15244_ _15244_/A _15244_/B vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_110_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18398_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ hold5709/X _11789_/B _11406_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ hold799/X _15179_/B vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or2_1
X_12387_ hold35/X hold594/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14126_ _15525_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__or2_1
X_11338_ hold4911/X _12299_/B _11337_/X _12666_/A vssd1 vssd1 vccd1 vccd1 _11338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ hold1288/X _14105_/A2 _14056_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 _14057_/X
+ sky130_fd_sc_hd__o211a_1
X_11269_ hold4107/X _11747_/B _11268_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13008_ hold1467/X _13003_/Y _13007_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13008_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ _17877_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_1
X_17747_ _17747_/CLK _17747_/D vssd1 vssd1 vccd1 vccd1 _17747_/Q sky130_fd_sc_hd__dfxtp_1
X_14959_ hold2118/X _14946_/B _14958_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ _15539_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08480_/X sky130_fd_sc_hd__or2_1
X_17678_ _17678_/CLK _17678_/D vssd1 vssd1 vccd1 vccd1 _17678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16629_ _18233_/CLK _16629_/D vssd1 vssd1 vccd1 vccd1 _16629_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_269_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ hold2250/X _09106_/B _09100_/Y _14364_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09032_ hold214/X hold391/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__clkbuf_2
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 input46/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold344 hold344/A vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 hold366/A vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 hold377/A vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 hold388/A vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout802 fanout816/X vssd1 vssd1 vccd1 vccd1 _15003_/C1 sky130_fd_sc_hd__buf_4
X_09934_ hold5377/X _10028_/B _09933_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09934_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 _14939_/C1 vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__buf_4
Xfanout824 _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__buf_4
Xfanout835 _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14887_/C1 sky130_fd_sc_hd__buf_4
Xfanout846 _11791_/A vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__buf_6
X_09865_ hold4309/X _10049_/B _09864_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09865_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout857 _13312_/B1 vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__buf_6
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 input37/X vssd1 vssd1 vccd1 vccd1 hold943/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 _14950_/A vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__buf_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _08398_/X vssd1 vssd1 vccd1 vccd1 _15829_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 _15199_/A vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__buf_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _15751_/Q vssd1 vssd1 vccd1 vccd1 hold1022/X sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ hold26/X hold537/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__mux2_1
Xhold1033 _08389_/X vssd1 vssd1 vccd1 vccd1 _15826_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 _14173_/X vssd1 vssd1 vccd1 vccd1 _17889_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ hold5528/X _10780_/A2 _09795_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _09796_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _14412_/X vssd1 vssd1 vccd1 vccd1 _18004_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _13979_/X vssd1 vssd1 vccd1 vccd1 _17796_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ hold126/X hold424/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__mux2_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _17863_/Q vssd1 vssd1 vccd1 vccd1 hold1077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _17756_/Q vssd1 vssd1 vccd1 vccd1 hold1088/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1099 _08419_/X vssd1 vssd1 vccd1 vccd1 hold1099/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _09021_/A hold316/X vssd1 vssd1 vccd1 vccd1 _15960_/D sky130_fd_sc_hd__and2_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _16704_/Q _10640_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__and3_1
XFILLER_0_193_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _16681_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _13822_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_107_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ _17587_/Q _17121_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ hold4669/X _12341_/B _12240_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ hold4718/X _12356_/B _12171_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12172_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11123_ hold743/X hold4363/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__mux2_1
X_16980_ _17862_/CLK _16980_/D vssd1 vssd1 vccd1 vccd1 _16980_/Q sky130_fd_sc_hd__dfxtp_1
X_15931_ _17323_/CLK _15931_/D vssd1 vssd1 vccd1 vccd1 hold643/A sky130_fd_sc_hd__dfxtp_1
X_11054_ hold1124/X hold3940/X _11156_/C vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__mux2_1
X_10005_ _13126_/A _09933_/A _10004_/X vssd1 vssd1 vccd1 vccd1 _10005_/Y sky130_fd_sc_hd__a21oi_1
X_15862_ _17739_/CLK _15862_/D vssd1 vssd1 vccd1 vccd1 _15862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2290 _16250_/Q vssd1 vssd1 vccd1 vccd1 hold2290/X sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _17697_/CLK _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14813_ hold2776/X _14828_/B _14812_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14813_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _17692_/CLK _15793_/D vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17532_ _18308_/CLK _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_1
X_14744_ _15191_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__or2_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ hold5397/X _12338_/B _11955_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11956_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17463_ _17464_/CLK _17463_/D vssd1 vssd1 vccd1 vccd1 _17463_/Q sky130_fd_sc_hd__dfxtp_1
X_10907_ hold2913/X hold4716/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__mux2_1
X_14675_ hold2499/X _14666_/B _14674_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14675_/X
+ sky130_fd_sc_hd__o211a_1
X_11887_ hold3370/X _12374_/B _11886_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ _18385_/CLK _16414_/D vssd1 vssd1 vccd1 vccd1 _16414_/Q sky130_fd_sc_hd__dfxtp_1
X_13626_ _13800_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ hold2920/X _16770_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__mux2_1
X_17394_ _18448_/CLK _17394_/D vssd1 vssd1 vccd1 vccd1 _17394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16345_ _18358_/CLK _16345_/D vssd1 vssd1 vccd1 vccd1 _16345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ _13779_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__or2_1
X_10769_ hold2801/X hold5617/X _11066_/S vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ _17347_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__or2_1
X_13488_ _13776_/A _13488_/B vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__or2_1
X_16276_ _17480_/CLK hold781/X vssd1 vssd1 vccd1 vccd1 _16276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18015_ _18461_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
X_15227_ _15227_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15227_/X sky130_fd_sc_hd__or2_1
X_12439_ hold380/X hold662/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12440_/B sky130_fd_sc_hd__mux2_1
Xhold4609 _16619_/Q vssd1 vssd1 vccd1 vccd1 hold4609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ hold1063/X _15161_/B _15157_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _15158_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3908 _13803_/Y vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3919 _17577_/Q vssd1 vssd1 vccd1 vccd1 hold3919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ hold585/X hold272/X vssd1 vssd1 vccd1 vccd1 _14138_/B sky130_fd_sc_hd__or2_4
X_15089_ _15197_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__or2_1
X_07980_ _15549_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ hold867/X _16374_/Q _10571_/C vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__mux2_1
X_08601_ hold68/X hold697/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ hold861/X _13278_/A _10481_/S vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__mux2_1
X_08532_ hold23/X hold322/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_188_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08463_ hold2795/X _08488_/B _08462_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _08463_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08394_ _08504_/A _15508_/A vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__or2_4
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09015_ _09021_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _16124_/D sky130_fd_sc_hd__and2_1
Xhold5800 output79/X vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5811 output73/X vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_12
Xhold5822 _17519_/Q vssd1 vssd1 vccd1 vccd1 hold5822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5833 _18414_/Q vssd1 vssd1 vccd1 vccd1 hold5833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5844 _16281_/Q vssd1 vssd1 vccd1 vccd1 hold5844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5855 hold5855/A vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5866 hold5945/X vssd1 vssd1 vccd1 vccd1 hold5866/X sky130_fd_sc_hd__buf_2
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5877 hold5877/A vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_12
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5888 _16931_/Q vssd1 vssd1 vccd1 vccd1 hold5888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5899 _16529_/Q vssd1 vssd1 vccd1 vccd1 hold5899/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _15485_/B1 vssd1 vssd1 vccd1 vccd1 _09362_/D sky130_fd_sc_hd__clkbuf_8
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__buf_8
Xfanout621 _09351_/Y vssd1 vssd1 vccd1 vccd1 _15486_/A2 sky130_fd_sc_hd__buf_6
Xfanout632 _08598_/B vssd1 vssd1 vccd1 vccd1 _12509_/A2 sky130_fd_sc_hd__clkbuf_8
X_09917_ _18376_/Q _16463_/Q _10028_/C vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__mux2_1
Xfanout643 fanout660/X vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__buf_4
XFILLER_0_186_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout654 _12666_/A vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__buf_4
Xfanout665 _08159_/A vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__buf_4
Xfanout676 _14147_/C1 vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__buf_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 fanout842/X vssd1 vssd1 vccd1 vccd1 _14418_/C1 sky130_fd_sc_hd__clkbuf_4
X_09848_ hold2981/X _16440_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__mux2_1
Xfanout698 _08585_/A vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ hold1567/X _16417_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__mux2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ hold2475/X _17094_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ hold1361/X _17441_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ _17071_/Q _11741_/B _11741_/C vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__and3_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ hold2824/X _17048_/Q _11672_/S vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__mux2_1
X_14460_ hold2985/X _14481_/B _14459_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14460_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10623_ hold3745/X _10527_/A _10622_/X vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__a21oi_1
X_13411_ hold4801/X _12311_/B _13410_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _13411_/X
+ sky130_fd_sc_hd__o211a_1
X_14391_ _14786_/A hold1989/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _17345_/CLK _16130_/D vssd1 vssd1 vccd1 vccd1 hold591/A sky130_fd_sc_hd__dfxtp_1
X_13342_ hold3997/X _13829_/B _13341_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10554_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _13273_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13273_/X sky130_fd_sc_hd__and2_1
X_16061_ _18408_/CLK _16061_/D vssd1 vssd1 vccd1 vccd1 hold448/A sky130_fd_sc_hd__dfxtp_1
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__or2_1
Xclkbuf_5_11__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_84_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_15012_ _15227_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__or2_1
X_12224_ hold1675/X _17232_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__mux2_1
X_12155_ hold2674/X hold4917/X _13388_/S vssd1 vssd1 vccd1 vccd1 _12156_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11106_/X sky130_fd_sc_hd__or2_1
X_12086_ hold2789/X _17186_/Q _13844_/C vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__mux2_1
X_16963_ _17907_/CLK _16963_/D vssd1 vssd1 vccd1 vccd1 _16963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15914_ _17289_/CLK _15914_/D vssd1 vssd1 vccd1 vccd1 hold390/A sky130_fd_sc_hd__dfxtp_1
X_11037_ _11067_/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11037_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16894_ _18065_/CLK _16894_/D vssd1 vssd1 vccd1 vccd1 _16894_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _17738_/CLK _15845_/D vssd1 vssd1 vccd1 vccd1 _15845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _17734_/CLK _15776_/D vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ hold1507/X _17507_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17516_/CLK _17515_/D vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_1
X_14727_ hold1836/X _14718_/B _14726_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14727_/X
+ sky130_fd_sc_hd__o211a_1
X_11939_ hold2528/X hold4569/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__mux2_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17446_ _17691_/CLK _17446_/D vssd1 vssd1 vccd1 vccd1 _17446_/Q sky130_fd_sc_hd__dfxtp_1
X_14658_ _15105_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13609_ hold4049/X _13805_/B _13608_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__o211a_1
X_17377_ _17480_/CLK _17377_/D vssd1 vssd1 vccd1 vccd1 _17377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ hold1597/X _14610_/B _14588_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14589_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _18241_/CLK _16328_/D vssd1 vssd1 vccd1 vccd1 _16328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5107 _11881_/X vssd1 vssd1 vccd1 vccd1 _17117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5118 _16513_/Q vssd1 vssd1 vccd1 vccd1 hold5118/X sky130_fd_sc_hd__dlygate4sd3_1
X_16259_ _17485_/CLK _16259_/D vssd1 vssd1 vccd1 vccd1 _16259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5129 _11839_/X vssd1 vssd1 vccd1 vccd1 _17103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4406 _10921_/X vssd1 vssd1 vccd1 vccd1 _16797_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4417 _17661_/Q vssd1 vssd1 vccd1 vccd1 hold4417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4428 _12289_/X vssd1 vssd1 vccd1 vccd1 _17253_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4439 _17212_/Q vssd1 vssd1 vccd1 vccd1 hold4439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3705 _16737_/Q vssd1 vssd1 vccd1 vccd1 hold3705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3716 _16349_/Q vssd1 vssd1 vccd1 vccd1 _13262_/A sky130_fd_sc_hd__buf_1
Xhold3727 _10033_/Y vssd1 vssd1 vccd1 vccd1 _16501_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3738 _11730_/Y vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3749 _10593_/Y vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07963_ hold1251/X _07978_/B _07962_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _07963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09702_ _09903_/A _09702_/B vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07894_ _14511_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09633_ _10779_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_284_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17908_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09564_ _09954_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_213_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18025_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08515_ _15519_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _14555_/B _14555_/C _09495_/C vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__or3_1
XFILLER_0_78_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ hold2020/X _08433_/B _08445_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _08379_/A hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__and2_1
XFILLER_0_147_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5630 _10912_/X vssd1 vssd1 vccd1 vccd1 _16794_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5641 _16425_/Q vssd1 vssd1 vccd1 vccd1 hold5641/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ hold4297/X _11192_/B _10269_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10270_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5652 _11125_/X vssd1 vssd1 vccd1 vccd1 _16865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5663 _11032_/X vssd1 vssd1 vccd1 vccd1 _16834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5674 _16898_/Q vssd1 vssd1 vccd1 vccd1 hold5674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4940 _11413_/X vssd1 vssd1 vccd1 vccd1 _16961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5685 _16867_/Q vssd1 vssd1 vccd1 vccd1 hold5685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4951 _17261_/Q vssd1 vssd1 vccd1 vccd1 hold4951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5696 _09598_/X vssd1 vssd1 vccd1 vccd1 _16356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4962 _12262_/X vssd1 vssd1 vccd1 vccd1 _17244_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4973 _17275_/Q vssd1 vssd1 vccd1 vccd1 hold4973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4984 _13741_/X vssd1 vssd1 vccd1 vccd1 _17700_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4995 _17724_/Q vssd1 vssd1 vccd1 vccd1 hold4995/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout440 fanout484/X vssd1 vssd1 vccd1 vccd1 _12308_/C sky130_fd_sc_hd__buf_4
Xfanout451 fanout484/X vssd1 vssd1 vccd1 vccd1 _11717_/C sky130_fd_sc_hd__buf_4
Xfanout462 _12332_/C vssd1 vssd1 vccd1 vccd1 _13871_/C sky130_fd_sc_hd__clkbuf_8
Xfanout473 _11672_/S vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__buf_4
X_13960_ _15521_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13960_/X sky130_fd_sc_hd__or2_1
Xfanout484 _09499_/Y vssd1 vssd1 vccd1 vccd1 fanout484/X sky130_fd_sc_hd__buf_8
Xfanout495 _10001_/C vssd1 vssd1 vccd1 vccd1 _10025_/C sky130_fd_sc_hd__clkbuf_8
X_12911_ hold3006/X _12910_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__mux2_1
X_13891_ hold241/X hold271/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__nor2_1
X_15630_ _18445_/CLK _15630_/D vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ hold3080/X _12841_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__mux2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _17718_/CLK _15561_/D vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12773_ hold3458/X _12772_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__mux2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17300_/CLK _17300_/D vssd1 vssd1 vccd1 vccd1 hold395/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ hold971/X _14554_/A2 _14511_/X _13901_/A vssd1 vssd1 vccd1 vccd1 hold972/A
+ sky130_fd_sc_hd__o211a_1
X_18280_ _18416_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ hold3787/X _11631_/A _11723_/X vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15492_/A hold242/X vssd1 vssd1 vccd1 vccd1 _15505_/S sky130_fd_sc_hd__nand2_8
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17231_ _17263_/CLK _17231_/D vssd1 vssd1 vccd1 vccd1 _17231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _12234_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
X_14443_ _15231_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17345_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10606_ _10651_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10606_/Y sky130_fd_sc_hd__nor2_1
X_17162_ _18445_/CLK _17162_/D vssd1 vssd1 vccd1 vccd1 _17162_/Q sky130_fd_sc_hd__dfxtp_1
X_11586_ _12093_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__or2_1
X_14374_ _15036_/A _14374_/B vssd1 vssd1 vccd1 vccd1 _17986_/D sky130_fd_sc_hd__and2_1
XFILLER_0_141_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ _18409_/CLK _16113_/D vssd1 vssd1 vccd1 vccd1 hold361/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10537_ hold4571/X _10631_/B _10536_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10537_/X
+ sky130_fd_sc_hd__o211a_1
X_13325_ hold1302/X hold3865/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17093_ _17253_/CLK _17093_/D vssd1 vssd1 vccd1 vccd1 _17093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _18423_/CLK _16044_/D vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
X_13256_ _13249_/X _13255_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__o21a_1
X_10468_ hold3531/X _11192_/B _10467_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _13716_/A _12207_/B vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__or2_1
X_13187_ _13186_/X _16916_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__mux2_1
X_10399_ hold4157/X _10589_/B _10398_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10399_/X
+ sky130_fd_sc_hd__o211a_1
X_12138_ _12234_/A _12138_/B vssd1 vssd1 vccd1 vccd1 _12138_/X sky130_fd_sc_hd__or2_1
X_17995_ _18061_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
X_12069_ _13392_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
X_16946_ _17889_/CLK _16946_/D vssd1 vssd1 vccd1 vccd1 _16946_/Q sky130_fd_sc_hd__dfxtp_1
X_16877_ _18071_/CLK _16877_/D vssd1 vssd1 vccd1 vccd1 _16877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _17719_/CLK _15828_/D vssd1 vssd1 vccd1 vccd1 _15828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15759_ _17678_/CLK _15759_/D vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfxtp_1
X_08300_ hold1027/X _08336_/A2 _08299_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _08300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09280_ _12813_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _16251_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ hold1227/X _08262_/B _08230_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17429_ _17691_/CLK _17429_/D vssd1 vssd1 vccd1 vccd1 _17429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _15513_/A hold2475/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ hold1455/X _08088_/B _08092_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4203 _16600_/Q vssd1 vssd1 vccd1 vccd1 hold4203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4214 _10402_/X vssd1 vssd1 vccd1 vccd1 _16624_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4225 _10168_/X vssd1 vssd1 vccd1 vccd1 _16546_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4236 _16667_/Q vssd1 vssd1 vccd1 vccd1 hold4236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3502 _16649_/Q vssd1 vssd1 vccd1 vccd1 hold3502/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4247 _10120_/X vssd1 vssd1 vccd1 vccd1 _16530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3513 _17685_/Q vssd1 vssd1 vccd1 vccd1 hold3513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4258 _10846_/X vssd1 vssd1 vccd1 vccd1 _16772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3524 _16555_/Q vssd1 vssd1 vccd1 vccd1 hold3524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4269 _17038_/Q vssd1 vssd1 vccd1 vccd1 hold4269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3535 _16415_/Q vssd1 vssd1 vccd1 vccd1 hold3535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3546 _17447_/Q vssd1 vssd1 vccd1 vccd1 hold3546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2801 _17950_/Q vssd1 vssd1 vccd1 vccd1 hold2801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 _08298_/X vssd1 vssd1 vccd1 vccd1 _15782_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3557 _13582_/X vssd1 vssd1 vccd1 vccd1 _17647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ hold14/X hold528/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__mux2_1
Xhold3568 _17745_/Q vssd1 vssd1 vccd1 vccd1 _13874_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2823 _14420_/X vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2834 _17883_/Q vssd1 vssd1 vccd1 vccd1 hold2834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3579 _17671_/Q vssd1 vssd1 vccd1 vccd1 hold3579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2845 _14257_/X vssd1 vssd1 vccd1 vccd1 _17929_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2856 _18334_/Q vssd1 vssd1 vccd1 vccd1 hold2856/X sky130_fd_sc_hd__dlygate4sd3_1
X_07946_ _14850_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07946_/X sky130_fd_sc_hd__or2_1
Xhold2867 _14510_/X vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2878 _18024_/Q vssd1 vssd1 vccd1 vccd1 hold2878/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2889 _18034_/Q vssd1 vssd1 vccd1 vccd1 hold2889/X sky130_fd_sc_hd__dlygate4sd3_1
X_07877_ hold800/X _07881_/B vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__or2_1
X_09616_ hold5647/X _09992_/B _09615_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09616_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ hold5498/X _10025_/B _09546_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09547_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09478_ _09483_/C _09481_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _16320_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08429_ _15217_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ hold4205/X _11726_/B _11439_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11371_ hold5580/X _11753_/B _11370_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11371_/X
+ sky130_fd_sc_hd__o211a_1
X_13110_ _13110_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__or2_1
X_10322_ hold2409/X _16598_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__mux2_1
X_14090_ _15543_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _17522_/Q hold793/X _17523_/Q vssd1 vssd1 vccd1 vccd1 hold794/A sky130_fd_sc_hd__or3b_1
Xhold5460 _17010_/Q vssd1 vssd1 vccd1 vccd1 hold5460/X sky130_fd_sc_hd__dlygate4sd3_1
X_10253_ hold2685/X _16575_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__mux2_1
Xhold5471 _11662_/X vssd1 vssd1 vccd1 vccd1 _17044_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5482 _16403_/Q vssd1 vssd1 vccd1 vccd1 hold5482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5493 _09766_/X vssd1 vssd1 vccd1 vccd1 _16412_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4770 _11821_/X vssd1 vssd1 vccd1 vccd1 _17097_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10184_ hold2973/X _16552_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__mux2_1
Xhold4781 _17233_/Q vssd1 vssd1 vccd1 vccd1 hold4781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4792 _10804_/X vssd1 vssd1 vccd1 vccd1 _16758_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16800_ _18035_/CLK _16800_/D vssd1 vssd1 vccd1 vccd1 _16800_/Q sky130_fd_sc_hd__dfxtp_1
X_17780_ _18427_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_135_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18358_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14992_ _15207_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__or2_1
Xfanout270 _11076_/A vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__buf_4
Xfanout281 _13779_/A vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__buf_4
Xfanout292 _11697_/A vssd1 vssd1 vccd1 vccd1 _12153_/A sky130_fd_sc_hd__clkbuf_4
X_16731_ _18054_/CLK _16731_/D vssd1 vssd1 vccd1 vccd1 _16731_/Q sky130_fd_sc_hd__dfxtp_1
X_13943_ _13943_/A _13943_/B vssd1 vssd1 vccd1 vccd1 _17779_/D sky130_fd_sc_hd__and2_1
XFILLER_0_191_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ _18220_/CLK _16662_/D vssd1 vssd1 vccd1 vccd1 _16662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13874_ _13874_/A _13886_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13874_/X sky130_fd_sc_hd__and3_1
X_18401_ _18417_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
X_15613_ _17583_/CLK _15613_/D vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ _12825_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _17451_/D sky130_fd_sc_hd__and2_1
X_16593_ _18215_/CLK _16593_/D vssd1 vssd1 vccd1 vccd1 _16593_/Q sky130_fd_sc_hd__dfxtp_1
X_18332_ _18388_/CLK hold938/X vssd1 vssd1 vccd1 vccd1 hold937/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ hold1985/X _15547_/B _15543_/Y _12666_/A vssd1 vssd1 vccd1 vccd1 _15544_/X
+ sky130_fd_sc_hd__o211a_1
X_12756_ _12756_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _17428_/D sky130_fd_sc_hd__and2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ hold4929/X _12341_/B _11706_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11707_/X
+ sky130_fd_sc_hd__o211a_1
X_18263_ _18385_/CLK hold848/X vssd1 vssd1 vccd1 vccd1 hold847/A sky130_fd_sc_hd__dfxtp_1
X_15475_ hold580/X _09386_/A _09362_/D hold525/X vssd1 vssd1 vccd1 vccd1 _15475_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ _12789_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _17405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17214_ _17266_/CLK _17214_/D vssd1 vssd1 vccd1 vccd1 _17214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14426_ hold1306/X _14433_/B _14425_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _14426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18194_ _18226_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11638_ hold4887/X _11732_/B _11637_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11638_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _17583_/CLK _17145_/D vssd1 vssd1 vccd1 vccd1 _17145_/Q sky130_fd_sc_hd__dfxtp_1
X_14357_ _14984_/A hold2729/X hold275/X vssd1 vssd1 vccd1 vccd1 _14358_/B sky130_fd_sc_hd__mux2_1
X_11569_ hold4121/X _11798_/B _11568_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold707 hold707/A vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 hold718/A vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ hold5300/X _13307_/X _13308_/S vssd1 vssd1 vccd1 vccd1 _13308_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold729 hold740/X vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ _17862_/CLK _17076_/D vssd1 vssd1 vccd1 vccd1 _17076_/Q sky130_fd_sc_hd__dfxtp_1
X_14288_ _15183_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14288_/X sky130_fd_sc_hd__or2_1
X_16027_ _18425_/CLK _16027_/D vssd1 vssd1 vccd1 vccd1 hold537/A sky130_fd_sc_hd__dfxtp_1
X_13239_ _13311_/A1 _13237_/X _13238_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2108 _15827_/Q vssd1 vssd1 vccd1 vccd1 hold2108/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 _14959_/X vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07800_ _18461_/Q _18459_/Q vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__nor2_1
X_08780_ _15414_/A hold252/X vssd1 vssd1 vccd1 vccd1 _16010_/D sky130_fd_sc_hd__and2_1
Xhold1407 _16249_/Q vssd1 vssd1 vccd1 vccd1 hold1407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _15757_/Q vssd1 vssd1 vccd1 vccd1 hold1418/X sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ _18431_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1429 _13991_/X vssd1 vssd1 vccd1 vccd1 _17802_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16929_ _17777_/CLK _16929_/D vssd1 vssd1 vccd1 vccd1 _16929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _15231_/A _07804_/B _09401_/S vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09332_ hold5981/X _09338_/A2 hold780/X _12909_/A vssd1 vssd1 vccd1 vccd1 hold781/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _15539_/A hold917/X _09277_/S vssd1 vssd1 vccd1 vccd1 hold918/A sky130_fd_sc_hd__mux2_1
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08214_ hold2216/X _08213_/B _08213_/Y _08257_/C1 vssd1 vssd1 vccd1 vccd1 _08214_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ hold949/X _09228_/B vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ _08147_/A _08145_/B vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08076_ _14529_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4000 _09619_/X vssd1 vssd1 vccd1 vccd1 _16363_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4011 _10786_/X vssd1 vssd1 vccd1 vccd1 _16752_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4022 _16690_/Q vssd1 vssd1 vccd1 vccd1 hold4022/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4033 _16577_/Q vssd1 vssd1 vccd1 vccd1 hold4033/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4044 _11062_/X vssd1 vssd1 vccd1 vccd1 _16844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4055 _17729_/Q vssd1 vssd1 vccd1 vccd1 hold4055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3310 _12860_/X vssd1 vssd1 vccd1 vccd1 _12861_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4066 _10555_/X vssd1 vssd1 vccd1 vccd1 _16675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3321 _11824_/X vssd1 vssd1 vccd1 vccd1 _17098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3332 _17255_/Q vssd1 vssd1 vccd1 vccd1 hold3332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4077 _16822_/Q vssd1 vssd1 vccd1 vccd1 hold4077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3343 _10237_/X vssd1 vssd1 vccd1 vccd1 _16569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4088 _11356_/X vssd1 vssd1 vccd1 vccd1 _16942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3354 _11932_/X vssd1 vssd1 vccd1 vccd1 _17134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4099 _17054_/Q vssd1 vssd1 vccd1 vccd1 hold4099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3365 _10525_/X vssd1 vssd1 vccd1 vccd1 _16665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2620 _17815_/Q vssd1 vssd1 vccd1 vccd1 hold2620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__buf_4
Xhold2631 _17908_/Q vssd1 vssd1 vccd1 vccd1 hold2631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3376 _17048_/Q vssd1 vssd1 vccd1 vccd1 hold3376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3387 _09565_/X vssd1 vssd1 vccd1 vccd1 _16345_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2642 _14540_/X vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _15414_/A hold102/X vssd1 vssd1 vccd1 vccd1 _16106_/D sky130_fd_sc_hd__and2_1
Xhold2653 _09227_/X vssd1 vssd1 vccd1 vccd1 _16225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3398 _16416_/Q vssd1 vssd1 vccd1 vccd1 hold3398/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__clkbuf_2
Xhold2664 _17946_/Q vssd1 vssd1 vccd1 vccd1 hold2664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1930 _15685_/Q vssd1 vssd1 vccd1 vccd1 hold1930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 _07899_/X vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__clkbuf_2
Xhold2686 _14683_/X vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ hold1519/X _07924_/B _07928_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _07929_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1941 _17829_/Q vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1952 _18153_/Q vssd1 vssd1 vccd1 vccd1 hold1952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2697 _16172_/Q vssd1 vssd1 vccd1 vccd1 hold2697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 _15168_/X vssd1 vssd1 vccd1 vccd1 _18367_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _14661_/X vssd1 vssd1 vccd1 vccd1 _18123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1985 _18450_/Q vssd1 vssd1 vccd1 vccd1 hold1985/X sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ _18007_/Q _16804_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__mux2_1
Xhold1996 _18184_/Q vssd1 vssd1 vccd1 vccd1 hold1996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ hold2167/X _16781_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ hold2151/X hold3124/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13791_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__or2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ hold2644/X _17358_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15260_ hold164/X _15486_/A2 _15446_/B1 hold454/X vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _17329_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ hold2631/X _14198_/B _14210_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14211_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11423_ hold2658/X _16965_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__mux2_1
X_15191_ _15191_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _13132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14142_ _15000_/A hold587/X vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__nand2_1
X_11354_ hold2417/X hold4020/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11355_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _10563_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14073_ hold1253/X _14105_/A2 _14072_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _14073_/X
+ sky130_fd_sc_hd__o211a_1
X_11285_ hold1319/X hold5331/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_316_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17721_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5290 _11776_/Y vssd1 vssd1 vccd1 vccd1 _17082_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13024_ _17518_/Q hold901/X vssd1 vssd1 vccd1 vccd1 hold902/A sky130_fd_sc_hd__nand2_1
X_10236_ _10422_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__or2_1
X_17901_ _17901_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_1
X_17832_ _17896_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
X_10167_ _10521_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__or2_1
X_17763_ _17827_/CLK _17763_/D vssd1 vssd1 vccd1 vccd1 _17763_/Q sky130_fd_sc_hd__dfxtp_1
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__or2_1
X_14975_ hold685/X _15006_/B _14974_/X _15044_/A vssd1 vssd1 vccd1 vccd1 hold686/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16714_ _18042_/CLK _16714_/D vssd1 vssd1 vccd1 vccd1 _16714_/Q sky130_fd_sc_hd__dfxtp_1
X_13926_ hold265/A _17771_/Q hold244/X vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__mux2_1
X_17694_ _17694_/CLK _17694_/D vssd1 vssd1 vccd1 vccd1 _17694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16645_ _18235_/CLK _16645_/D vssd1 vssd1 vccd1 vccd1 _16645_/Q sky130_fd_sc_hd__dfxtp_1
X_13857_ hold3770/X _13764_/A _13856_/X vssd1 vssd1 vccd1 vccd1 _13857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12808_ hold1710/X _17447_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux2_1
X_16576_ _18198_/CLK _16576_/D vssd1 vssd1 vccd1 vccd1 _16576_/Q sky130_fd_sc_hd__dfxtp_1
X_13788_ _13788_/A _13788_/B vssd1 vssd1 vccd1 vccd1 _13788_/X sky130_fd_sc_hd__or2_1
X_18315_ _18315_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__dfxtp_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _15527_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15527_/X sky130_fd_sc_hd__or2_1
X_12739_ _16244_/Q hold3035/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18043_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18246_ _18420_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
X_15458_ hold643/X _09367_/A _09362_/C hold644/X vssd1 vssd1 vccd1 vccd1 _15458_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ _14517_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__or2_1
X_18177_ _18268_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ hold132/X _09365_/B _09392_/C hold507/X _15388_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _17128_/CLK _17128_/D vssd1 vssd1 vccd1 vccd1 _17128_/Q sky130_fd_sc_hd__dfxtp_1
Xhold515 hold515/A vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold526 hold526/A vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold537 hold537/A vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 hold548/A vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ hold1768/X hold5072/X _10271_/S vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__mux2_1
Xhold559 hold559/A vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _17907_/CLK _17059_/D vssd1 vssd1 vccd1 vccd1 _17059_/Q sky130_fd_sc_hd__dfxtp_1
X_08901_ _15374_/A _08901_/B vssd1 vssd1 vccd1 vccd1 _16068_/D sky130_fd_sc_hd__and2_1
X_09881_ hold1267/X hold5098/X _10481_/S vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ hold71/X hold648/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _17893_/Q vssd1 vssd1 vccd1 vccd1 hold1204/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _07949_/X vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _08467_/X vssd1 vssd1 vccd1 vccd1 _15862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _16156_/Q vssd1 vssd1 vccd1 vccd1 hold1237/X sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ hold214/X _16002_/Q _08787_/S vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__mux2_1
Xhold1248 _17981_/Q vssd1 vssd1 vccd1 vccd1 hold1248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 la_data_in[12] vssd1 vssd1 vccd1 vccd1 hold1259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _09003_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _15968_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _15103_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _12777_/A _09246_/B vssd1 vssd1 vccd1 vccd1 _16234_/D sky130_fd_sc_hd__and2_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ hold2121/X _09177_/A2 _09176_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08128_ _15533_/A hold2480/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ hold1497/X _08082_/B _08058_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _08059_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11070_ _11106_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__or2_1
Xoutput79 _13185_/A vssd1 vssd1 vccd1 vccd1 output79/X sky130_fd_sc_hd__buf_6
XFILLER_0_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3140 _13864_/Y vssd1 vssd1 vccd1 vccd1 _17741_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10021_ _11203_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10021_/Y sky130_fd_sc_hd__nor2_1
Xhold3151 _13809_/Y vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3162 _17119_/Q vssd1 vssd1 vccd1 vccd1 hold3162/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3173 _10069_/Y vssd1 vssd1 vccd1 vccd1 _16513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3184 _11719_/Y vssd1 vssd1 vccd1 vccd1 _17063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2450 _08008_/X vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3195 _10978_/X vssd1 vssd1 vccd1 vccd1 _16816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2461 _15808_/Q vssd1 vssd1 vccd1 vccd1 hold2461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2472 _08012_/X vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _16268_/Q vssd1 vssd1 vccd1 vccd1 hold2483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2494 _14069_/X vssd1 vssd1 vccd1 vccd1 _17839_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 _18446_/Q vssd1 vssd1 vccd1 vccd1 hold1760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1771 input1/X vssd1 vssd1 vccd1 vccd1 hold1771/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _15099_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__or2_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ hold1968/X hold4597/X _13871_/C vssd1 vssd1 vccd1 vccd1 _11973_/B sky130_fd_sc_hd__mux2_1
Xhold1782 _09314_/X vssd1 vssd1 vccd1 vccd1 _16267_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _07925_/X vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ hold4807/X _13805_/B _13710_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13711_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _11667_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__or2_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ hold1436/X _14718_/B _14690_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14691_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _18416_/CLK _16430_/D vssd1 vssd1 vccd1 vccd1 _16430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13642_ hold4345/X _13832_/B _13641_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13642_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10854_ _11616_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _18243_/CLK _16361_/D vssd1 vssd1 vccd1 vccd1 _16361_/Q sky130_fd_sc_hd__dfxtp_1
X_13573_ hold5173/X _13859_/B _13572_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13573_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _11652_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10785_/X sky130_fd_sc_hd__or2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _18222_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
X_15312_ _15471_/A _15312_/B _15312_/C _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/X
+ sky130_fd_sc_hd__or4_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ hold3465/X _12523_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__mux2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16314_/CLK _16292_/D vssd1 vssd1 vccd1 vccd1 _16292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _18063_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _15490_/A1 _15235_/X _15242_/X _15490_/B1 hold3989/X vssd1 vssd1 vccd1 vccd1
+ _15243_/X sky130_fd_sc_hd__a32o_1
X_12455_ hold32/X _08598_/B _08999_/B _12454_/X _15454_/A vssd1 vssd1 vccd1 vccd1
+ hold33/A sky130_fd_sc_hd__o311a_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ _11694_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15174_ hold853/X hold609/X _15173_/X _15394_/A vssd1 vssd1 vccd1 vccd1 hold854/A
+ sky130_fd_sc_hd__o211a_1
X_12386_ _15414_/A hold408/X vssd1 vssd1 vccd1 vccd1 _17286_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14125_ hold1309/X hold587/X _14124_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _14125_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11337_ _12204_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_150_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18183_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14056_ hold944/X _14072_/B vssd1 vssd1 vccd1 vccd1 _14056_/X sky130_fd_sc_hd__or2_1
X_11268_ _11652_/A _11268_/B vssd1 vssd1 vccd1 vccd1 _11268_/X sky130_fd_sc_hd__or2_1
X_13007_ _14970_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__or2_1
X_10219_ hold4516/X _10619_/B _10218_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _10219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ hold5297/X _11103_/A _11198_/X vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__a21oi_1
X_17815_ _17880_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17746_ _17749_/CLK _17746_/D vssd1 vssd1 vccd1 vccd1 _17746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _15227_/A _14962_/B vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__or2_1
X_13909_ _13909_/A _13909_/B vssd1 vssd1 vccd1 vccd1 _17762_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17677_ _17741_/CLK _17677_/D vssd1 vssd1 vccd1 vccd1 _17677_/Q sky130_fd_sc_hd__dfxtp_1
X_14889_ hold2016/X _14880_/B _14888_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/X
+ sky130_fd_sc_hd__o211a_1
X_16628_ _18218_/CLK _16628_/D vssd1 vssd1 vccd1 vccd1 _16628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ _18149_/CLK _16559_/D vssd1 vssd1 vccd1 vccd1 _16559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09100_ _15541_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ _15414_/A hold180/X vssd1 vssd1 vccd1 vccd1 _16132_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18229_ _18229_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_238_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17747_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__clkbuf_2
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold334 input46/X vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold345 hold440/X vssd1 vssd1 vccd1 vccd1 hold441/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 hold61/X vssd1 vssd1 vccd1 vccd1 input26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 hold389/A vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__or2_1
Xfanout803 _15066_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__buf_4
Xfanout814 _14939_/C1 vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__buf_4
Xfanout825 fanout841/X vssd1 vssd1 vccd1 vccd1 _14733_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout836 _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14883_/C1 sky130_fd_sc_hd__buf_4
X_09864_ _10098_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__or2_1
Xfanout847 _11791_/A vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__clkbuf_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 _13312_/B1 vssd1 vssd1 vccd1 vccd1 _13304_/B1 sky130_fd_sc_hd__clkbuf_8
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _14504_/X vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _14950_/A vssd1 vssd1 vccd1 vccd1 _15219_/A sky130_fd_sc_hd__clkbuf_16
Xhold1012 hold5837/X vssd1 vssd1 vccd1 vccd1 _13053_/A sky130_fd_sc_hd__buf_4
X_08815_ _12422_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _16026_/D sky130_fd_sc_hd__and2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _08233_/X vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 _18427_/Q vssd1 vssd1 vccd1 vccd1 hold1034/X sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _11106_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__or2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1045 la_data_in[9] vssd1 vssd1 vccd1 vccd1 hold881/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 hold1296/X vssd1 vssd1 vccd1 vccd1 hold1297/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _16254_/Q vssd1 vssd1 vccd1 vccd1 hold1067/X sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _15334_/A hold159/X vssd1 vssd1 vccd1 vccd1 _15993_/D sky130_fd_sc_hd__and2_1
Xhold1078 _14119_/X vssd1 vssd1 vccd1 vccd1 _17863_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _17511_/Q vssd1 vssd1 vccd1 vccd1 hold1089/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ hold26/X _15960_/Q _08721_/S vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__mux2_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _11194_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10570_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ hold2750/X _09216_/B _09228_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_5_10__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_77_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_12240_ _12246_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _13392_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11122_ hold5393/X _11216_/B _11121_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _11122_/X
+ sky130_fd_sc_hd__o211a_1
Xhold890 input48/X vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__buf_1
X_15930_ _17523_/CLK _15930_/D vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__dfxtp_1
X_11053_ hold3929/X _11150_/B _11052_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _11053_/X
+ sky130_fd_sc_hd__o211a_1
X_10004_ _16492_/Q _10013_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__and3_1
X_15861_ _17739_/CLK _15861_/D vssd1 vssd1 vccd1 vccd1 _15861_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2280 _08489_/X vssd1 vssd1 vccd1 vccd1 _15873_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17600_ _17728_/CLK _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2291 _15575_/Q vssd1 vssd1 vccd1 vccd1 hold2291/X sky130_fd_sc_hd__dlygate4sd3_1
X_14812_ _15205_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__or2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _17723_/CLK _15792_/D vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17531_/CLK _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1590 _15132_/X vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ hold2846/X _14772_/B _14742_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14743_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _12051_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17462_ _17464_/CLK _17462_/D vssd1 vssd1 vccd1 vccd1 _17462_/Q sky130_fd_sc_hd__dfxtp_1
X_10906_ hold5550/X _11213_/B _10905_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10906_/X
+ sky130_fd_sc_hd__o211a_1
X_14674_ _14728_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _12279_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__or2_1
X_16413_ _18390_/CLK _16413_/D vssd1 vssd1 vccd1 vccd1 _16413_/Q sky130_fd_sc_hd__dfxtp_1
X_13625_ hold1820/X _17662_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17393_ _18456_/CLK _17393_/D vssd1 vssd1 vccd1 vccd1 _17393_/Q sky130_fd_sc_hd__dfxtp_1
X_10837_ hold4353/X _11222_/B _10836_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _10837_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ _18176_/CLK _16344_/D vssd1 vssd1 vccd1 vccd1 _16344_/Q sky130_fd_sc_hd__dfxtp_1
X_13556_ hold1842/X hold3577/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ hold5445/X _11150_/B _10767_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ hold14/X _12509_/A2 _12445_/B _12506_/X _12420_/A vssd1 vssd1 vccd1 vccd1
+ hold15/A sky130_fd_sc_hd__o311a_1
XFILLER_0_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16275_ _17480_/CLK _16275_/D vssd1 vssd1 vccd1 vccd1 _16275_/Q sky130_fd_sc_hd__dfxtp_1
X_13487_ hold2020/X hold4589/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13488_/B sky130_fd_sc_hd__mux2_1
X_10699_ hold5084/X _11177_/B _10698_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18014_ _18046_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_29__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_29__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_15226_ hold1718/X _15221_/B _15225_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15226_/X
+ sky130_fd_sc_hd__o211a_1
X_12438_ _12438_/A _12438_/B vssd1 vssd1 vccd1 vccd1 _17312_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ hold735/X _15179_/B vssd1 vssd1 vccd1 vccd1 _15157_/X sky130_fd_sc_hd__or2_1
X_12369_ hold3147/X _12279_/A _12368_/X vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__a21oi_1
Xhold3909 _13804_/Y vssd1 vssd1 vccd1 vccd1 _17721_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14108_ hold585/X hold272/X vssd1 vssd1 vccd1 vccd1 hold586/A sky130_fd_sc_hd__nor2_1
X_15088_ hold1610/X _15113_/B _15087_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _15088_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ hold2197/X _14040_/B _14038_/Y _13901_/A vssd1 vssd1 vccd1 vccd1 _14039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08600_ _12402_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _15922_/D sky130_fd_sc_hd__and2_1
X_09580_ hold4307/X _10571_/B _09579_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09580_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08531_ _13046_/C _12380_/A vssd1 vssd1 vccd1 vccd1 _08562_/S sky130_fd_sc_hd__or2_2
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17729_ _17741_/CLK _17729_/D vssd1 vssd1 vccd1 vccd1 _17729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ _14246_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08393_ _08504_/A _15508_/A vssd1 vssd1 vccd1 vccd1 _08393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09014_ hold47/X hold294/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__mux2_1
Xhold5801 hold6037/X vssd1 vssd1 vccd1 vccd1 hold5801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5812 hold5933/X vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5823 _17520_/Q vssd1 vssd1 vccd1 vccd1 hold5823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5834 _18401_/Q vssd1 vssd1 vccd1 vccd1 hold5834/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold120 hold299/X vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__clkbuf_2
Xhold5845 hold5845/A vssd1 vssd1 vccd1 vccd1 hold5845/X sky130_fd_sc_hd__clkbuf_4
Xhold5856 _16285_/Q vssd1 vssd1 vccd1 vccd1 hold5856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5867 hold5867/A vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_12
Xhold142 hold170/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold49/X vssd1 vssd1 vccd1 vccd1 input22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5878 _17752_/Q vssd1 vssd1 vccd1 vccd1 hold5878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5889 _16928_/Q vssd1 vssd1 vccd1 vccd1 hold5889/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _12982_/S vssd1 vssd1 vccd1 vccd1 _13000_/S sky130_fd_sc_hd__clkbuf_8
Xfanout611 _09361_/Y vssd1 vssd1 vccd1 vccd1 _15485_/B1 sky130_fd_sc_hd__buf_6
X_09916_ hold5336/X _10028_/B _09915_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09916_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout622 _15485_/A2 vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__buf_6
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout633 _12445_/A vssd1 vssd1 vccd1 vccd1 _08598_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 _12831_/A vssd1 vssd1 vccd1 vccd1 _15534_/C1 sky130_fd_sc_hd__buf_4
Xfanout655 _12666_/A vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__buf_4
Xfanout666 _08159_/A vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__buf_4
X_09847_ hold4999/X _10049_/B _09846_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout677 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14147_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 _12951_/A vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__buf_4
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout699 _08585_/A vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ hold3446/X _10067_/B _09777_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09778_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _17519_/Q _17518_/Q vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__nand2b_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _12301_/A _11740_/B vssd1 vssd1 vccd1 vccd1 _11740_/Y sky130_fd_sc_hd__nor2_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ hold5705/X _11765_/B _11670_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11671_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13410_ _13794_/A _13410_/B vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10622_ _16698_/Q _10640_/B _10640_/C vssd1 vssd1 vccd1 vccd1 _10622_/X sky130_fd_sc_hd__and3_1
XFILLER_0_154_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14390_ _14390_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__and2_1
XFILLER_0_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13341_ _13734_/A _13341_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__or2_1
X_10553_ hold2016/X hold3221/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _18407_/CLK _16060_/D vssd1 vssd1 vccd1 vccd1 hold567/A sky130_fd_sc_hd__dfxtp_1
X_13272_ _13265_/X _13271_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__o21a_1
X_10484_ hold2266/X hold4079/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__mux2_1
X_15011_ hold1725/X _15004_/B _15010_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12223_ hold4824/X _12356_/B _12222_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ hold4862/X _13844_/B _12153_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _12154_/X
+ sky130_fd_sc_hd__o211a_1
X_11105_ hold2394/X hold5554/X _11201_/C vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__mux2_1
X_12085_ hold4869/X _12377_/B _12084_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12085_/X
+ sky130_fd_sc_hd__o211a_1
X_16962_ _17873_/CLK _16962_/D vssd1 vssd1 vccd1 vccd1 _16962_/Q sky130_fd_sc_hd__dfxtp_1
X_15913_ _17331_/CLK _15913_/D vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__dfxtp_1
X_11036_ hold1790/X hold3208/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11037_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16893_ _17798_/CLK _16893_/D vssd1 vssd1 vccd1 vccd1 _16893_/Q sky130_fd_sc_hd__dfxtp_1
X_15844_ _17735_/CLK _15844_/D vssd1 vssd1 vccd1 vccd1 _15844_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _17694_/CLK _15775_/D vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12987_/A _12987_/B vssd1 vssd1 vccd1 vccd1 _17505_/D sky130_fd_sc_hd__and2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14726_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__or2_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _17516_/CLK hold684/X vssd1 vssd1 vccd1 vccd1 hold683/A sky130_fd_sc_hd__dfxtp_1
X_11938_ hold4803/X _12320_/B _11937_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11938_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17445_ _17447_/CLK _17445_/D vssd1 vssd1 vccd1 vccd1 _17445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ hold2453/X _14664_/B _14656_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14657_/X
+ sky130_fd_sc_hd__o211a_1
X_11869_ hold4915/X _12347_/B _11868_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13608_ _13710_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _17480_/CLK _17376_/D vssd1 vssd1 vccd1 vccd1 _17376_/Q sky130_fd_sc_hd__dfxtp_1
X_14588_ _15197_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14588_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16327_ _18415_/CLK _16327_/D vssd1 vssd1 vccd1 vccd1 _16327_/Q sky130_fd_sc_hd__dfxtp_1
X_13539_ _13737_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _17379_/CLK _16258_/D vssd1 vssd1 vccd1 vccd1 _16258_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5108 _16825_/Q vssd1 vssd1 vccd1 vccd1 hold5108/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5119 _09973_/X vssd1 vssd1 vccd1 vccd1 _16481_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _15209_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4407 _16561_/Q vssd1 vssd1 vccd1 vccd1 hold4407/X sky130_fd_sc_hd__dlygate4sd3_1
X_16189_ _18432_/CLK _16189_/D vssd1 vssd1 vccd1 vccd1 _16189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4418 _13528_/X vssd1 vssd1 vccd1 vccd1 _17629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4429 _17009_/Q vssd1 vssd1 vccd1 vccd1 hold4429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3706 _11220_/Y vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3717 _10056_/Y vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3728 _16544_/Q vssd1 vssd1 vccd1 vccd1 hold3728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3739 _11731_/Y vssd1 vssd1 vccd1 vccd1 _17067_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07962_ _15531_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07962_/X sky130_fd_sc_hd__or2_1
X_09701_ hold2771/X hold5562/X _09998_/C vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__mux2_1
X_07893_ hold1694/X _07918_/B _07892_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _07893_/X
+ sky130_fd_sc_hd__o211a_1
X_09632_ hold2711/X _16368_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__mux2_1
X_09563_ hold831/X _16345_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ hold1302/X _08503_/Y _08513_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _08514_/X
+ sky130_fd_sc_hd__o211a_1
X_09494_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__or3_4
XFILLER_0_33_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ _14786_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_253_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17734_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08376_ hold335/A _15820_/Q hold122/X vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__mux2_1
XFILLER_0_163_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5620 _09964_/X vssd1 vssd1 vccd1 vccd1 _16478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5631 _16498_/Q vssd1 vssd1 vccd1 vccd1 hold5631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5642 _09709_/X vssd1 vssd1 vccd1 vccd1 _16393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5653 _17074_/Q vssd1 vssd1 vccd1 vccd1 hold5653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5664 _16485_/Q vssd1 vssd1 vccd1 vccd1 hold5664/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4930 _11707_/X vssd1 vssd1 vccd1 vccd1 _17059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5675 _11128_/X vssd1 vssd1 vccd1 vccd1 _16866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4941 _16995_/Q vssd1 vssd1 vccd1 vccd1 hold4941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5686 _11035_/X vssd1 vssd1 vccd1 vccd1 _16835_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4952 _12217_/X vssd1 vssd1 vccd1 vccd1 _17229_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5697 _16982_/Q vssd1 vssd1 vccd1 vccd1 hold5697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4963 _16963_/Q vssd1 vssd1 vccd1 vccd1 hold4963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4974 _12259_/X vssd1 vssd1 vccd1 vccd1 _17243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4985 _17200_/Q vssd1 vssd1 vccd1 vccd1 hold4985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4996 _13717_/X vssd1 vssd1 vccd1 vccd1 _17692_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout430 _13056_/X vssd1 vssd1 vccd1 vccd1 _13307_/S sky130_fd_sc_hd__buf_8
Xfanout441 _13862_/C vssd1 vssd1 vccd1 vccd1 _13829_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout452 _11741_/C vssd1 vssd1 vccd1 vccd1 _12320_/C sky130_fd_sc_hd__clkbuf_8
Xfanout463 _12332_/C vssd1 vssd1 vccd1 vccd1 _13388_/S sky130_fd_sc_hd__clkbuf_8
Xfanout474 _11210_/C vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__clkbuf_8
Xfanout485 _11156_/C vssd1 vssd1 vccd1 vccd1 _11153_/C sky130_fd_sc_hd__buf_6
Xfanout496 _10763_/S vssd1 vssd1 vccd1 vccd1 _10001_/C sky130_fd_sc_hd__buf_4
X_12910_ hold1381/X _17481_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
X_13890_ _14556_/A hold1119/X _09120_/Y hold928/X vssd1 vssd1 vccd1 vccd1 hold929/A
+ sky130_fd_sc_hd__a31o_1
X_12841_ hold2750/X hold3063/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__mux2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ hold2244/X _15560_/A2 _15559_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _15560_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ hold1101/X hold3455/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14511_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _17065_/Q _11726_/B _11726_/C vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__and3_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15491_ _15491_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17262_/CLK _17230_/D vssd1 vssd1 vccd1 vccd1 _17230_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ hold2361/X _14433_/B _14441_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ hold2909/X hold5504/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10605_ hold3132/X _10527_/A _10604_/X vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17161_ _17257_/CLK _17161_/D vssd1 vssd1 vccd1 vccd1 _17161_/Q sky130_fd_sc_hd__dfxtp_1
X_14373_ hold265/X hold399/X hold275/X vssd1 vssd1 vccd1 vccd1 _14374_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ hold2609/X hold4492/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16112_ _17523_/CLK _16112_/D vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__dfxtp_1
X_13324_ hold4897/X _13805_/B _13323_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__o211a_1
X_10536_ _10542_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17092_ _18426_/CLK _17092_/D vssd1 vssd1 vccd1 vccd1 _17092_/Q sky130_fd_sc_hd__dfxtp_1
X_16043_ _18414_/CLK _16043_/D vssd1 vssd1 vccd1 vccd1 hold507/A sky130_fd_sc_hd__dfxtp_1
X_13255_ _13311_/A1 _13253_/X _13254_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10557_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ hold2113/X hold4393/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__mux2_1
X_13186_ _17574_/Q _17108_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17516_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10398_ _10554_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12137_ hold1284/X hold5369/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__mux2_1
X_17994_ _18158_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12068_ hold1608/X _17180_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _12069_/B sky130_fd_sc_hd__mux2_1
X_16945_ _17889_/CLK _16945_/D vssd1 vssd1 vccd1 vccd1 _16945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11019_ _11667_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__or2_1
X_16876_ _18241_/CLK _16876_/D vssd1 vssd1 vccd1 vccd1 _16876_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _17715_/CLK _15827_/D vssd1 vssd1 vccd1 vccd1 _15827_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _17741_/CLK _15758_/D vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ hold1615/X _14718_/B _14708_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14709_/X
+ sky130_fd_sc_hd__o211a_1
X_15689_ _17744_/CLK _15689_/D vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08230_ hold944/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17428_ _17428_/CLK _17428_/D vssd1 vssd1 vccd1 vccd1 _17428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ _08161_/A hold893/X vssd1 vssd1 vccd1 vccd1 _15718_/D sky130_fd_sc_hd__and2_1
XFILLER_0_144_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17359_ _17379_/CLK _17359_/D vssd1 vssd1 vccd1 vccd1 _17359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08092_ _14330_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4204 _10234_/X vssd1 vssd1 vccd1 vccd1 _16568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4215 _17077_/Q vssd1 vssd1 vccd1 vccd1 _11759_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4226 _17693_/Q vssd1 vssd1 vccd1 vccd1 hold4226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4237 _10435_/X vssd1 vssd1 vccd1 vccd1 _16635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3503 _10381_/X vssd1 vssd1 vccd1 vccd1 _16617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4248 _16803_/Q vssd1 vssd1 vccd1 vccd1 hold4248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3514 _13600_/X vssd1 vssd1 vccd1 vccd1 _17653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4259 _17667_/Q vssd1 vssd1 vccd1 vccd1 hold4259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3525 _10099_/X vssd1 vssd1 vccd1 vccd1 _16523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3536 _09679_/X vssd1 vssd1 vccd1 vccd1 _16383_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2802 _14301_/X vssd1 vssd1 vccd1 vccd1 _17950_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08994_ _12402_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _16114_/D sky130_fd_sc_hd__and2_1
Xhold3547 _17432_/Q vssd1 vssd1 vccd1 vccd1 hold3547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2813 _15723_/Q vssd1 vssd1 vccd1 vccd1 hold2813/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3558 _16618_/Q vssd1 vssd1 vccd1 vccd1 hold3558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3569 _13780_/X vssd1 vssd1 vccd1 vccd1 _17713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 _17896_/Q vssd1 vssd1 vccd1 vccd1 hold2824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2835 _14159_/X vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2846 _18162_/Q vssd1 vssd1 vccd1 vccd1 hold2846/X sky130_fd_sc_hd__dlygate4sd3_1
X_07945_ hold2963/X _07991_/A2 _07944_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07945_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2857 _15100_/X vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2868 _18145_/Q vssd1 vssd1 vccd1 vccd1 hold2868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2879 _14454_/X vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07876_ hold1885/X _07869_/B _07875_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07876_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ _11067_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09924_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09477_/A hold681/X _09477_/C vssd1 vssd1 vccd1 vccd1 _09483_/C sky130_fd_sc_hd__and3_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ hold2425/X _08433_/B _08427_/Y _08389_/A vssd1 vssd1 vccd1 vccd1 _08428_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _15811_/D sky130_fd_sc_hd__and2_1
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11370_ _11658_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10321_ hold4051/X _10640_/B _10320_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5450 _16761_/Q vssd1 vssd1 vccd1 vccd1 hold5450/X sky130_fd_sc_hd__dlygate4sd3_1
X_13040_ input2/X input1/X hold792/X input3/X vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__or4b_1
Xhold5461 _11464_/X vssd1 vssd1 vccd1 vccd1 _16978_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10252_ hold4351/X _11213_/B _10251_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5472 _17235_/Q vssd1 vssd1 vccd1 vccd1 hold5472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5483 _09643_/X vssd1 vssd1 vccd1 vccd1 _16371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5494 _16958_/Q vssd1 vssd1 vccd1 vccd1 hold5494/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4760 _10309_/X vssd1 vssd1 vccd1 vccd1 _16593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10183_ hold5013/X _10568_/B _10182_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _10183_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4771 _16756_/Q vssd1 vssd1 vccd1 vccd1 hold4771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4782 _12133_/X vssd1 vssd1 vccd1 vccd1 _17201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4793 _17173_/Q vssd1 vssd1 vccd1 vccd1 hold4793/X sky130_fd_sc_hd__dlygate4sd3_1
X_14991_ hold2711/X _15006_/B _14990_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _14991_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout260 _12285_/A vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__buf_4
Xfanout271 _11076_/A vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__buf_4
Xfanout282 fanout298/X vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__clkbuf_4
X_13942_ _15123_/A _17779_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 _13942_/X sky130_fd_sc_hd__mux2_1
X_16730_ _18061_/CLK _16730_/D vssd1 vssd1 vccd1 vccd1 _16730_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout293 _11697_/A vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__buf_4
X_16661_ _18219_/CLK _16661_/D vssd1 vssd1 vccd1 vccd1 _16661_/Q sky130_fd_sc_hd__dfxtp_1
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _13873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_175_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18035_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18400_ _18409_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_15612_ _18426_/CLK _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfxtp_1
X_12824_ hold3083/X _12823_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__mux2_1
X_16592_ _18214_/CLK _16592_/D vssd1 vssd1 vccd1 vccd1 _16592_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17341_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18331_ _18395_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
X_15543_ _15543_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ hold3472/X _12754_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__mux2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18360_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _12246_/A _11706_/B vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__or2_1
X_15474_ _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__or2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ hold3092/X _12685_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _17743_/CLK _17213_/D vssd1 vssd1 vccd1 vccd1 _17213_/Q sky130_fd_sc_hd__dfxtp_1
X_14425_ _15105_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14425_/X sky130_fd_sc_hd__or2_1
X_18193_ _18225_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17144_ _17208_/CLK _17144_/D vssd1 vssd1 vccd1 vccd1 _17144_/Q sky130_fd_sc_hd__dfxtp_1
X_14356_ _14356_/A _14356_/B vssd1 vssd1 vccd1 vccd1 _17977_/D sky130_fd_sc_hd__and2_1
X_11568_ _12153_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__or2_1
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold708 hold708/A vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ _13306_/X hold5888/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__mux2_1
X_10519_ _10613_/A _10631_/B _10518_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10519_/X
+ sky130_fd_sc_hd__o211a_1
Xhold719 hold719/A vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ _17891_/CLK _17075_/D vssd1 vssd1 vccd1 vccd1 _17075_/Q sky130_fd_sc_hd__dfxtp_1
X_14287_ _15508_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14334_/B sky130_fd_sc_hd__or2_4
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _12234_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16026_ _17345_/CLK _16026_/D vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13238_ _13238_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13238_/X sky130_fd_sc_hd__or2_1
X_13169_ _13169_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__and2_1
XFILLER_0_62_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2109 _15580_/Q vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17977_ _18043_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1408 _18383_/Q vssd1 vssd1 vccd1 vccd1 hold1408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _08245_/X vssd1 vssd1 vccd1 vccd1 _15757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ _17893_/CLK _16928_/D vssd1 vssd1 vccd1 vccd1 _16928_/Q sky130_fd_sc_hd__dfxtp_1
X_16859_ _18054_/CLK _16859_/D vssd1 vssd1 vccd1 vccd1 _16859_/Q sky130_fd_sc_hd__dfxtp_1
X_09400_ _09400_/A hold801/X _09400_/C vssd1 vssd1 vccd1 vccd1 _09401_/S sky130_fd_sc_hd__or3_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ hold770/X _09337_/B vssd1 vssd1 vccd1 vccd1 hold780/A sky130_fd_sc_hd__or2_1
XFILLER_0_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _12756_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _16242_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08213_ _14774_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08213_/Y sky130_fd_sc_hd__nand2_1
X_09193_ hold2624/X _09216_/B _09192_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _09193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08144_ _15549_/A hold1876/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08145_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08075_ hold2528/X _08082_/B _08074_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _08075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4001 _16986_/Q vssd1 vssd1 vccd1 vccd1 hold4001/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4012 _16810_/Q vssd1 vssd1 vccd1 vccd1 hold4012/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4023 _10504_/X vssd1 vssd1 vccd1 vccd1 _16658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4034 _10165_/X vssd1 vssd1 vccd1 vccd1 _16545_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3300 _10981_/X vssd1 vssd1 vccd1 vccd1 _16817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4045 _16780_/Q vssd1 vssd1 vccd1 vccd1 hold4045/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3311 _16644_/Q vssd1 vssd1 vccd1 vccd1 hold3311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4056 _13732_/X vssd1 vssd1 vccd1 vccd1 _17697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3322 _17677_/Q vssd1 vssd1 vccd1 vccd1 hold3322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4067 _17663_/Q vssd1 vssd1 vccd1 vccd1 hold4067/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3333 _12199_/X vssd1 vssd1 vccd1 vccd1 _17223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4078 _10900_/X vssd1 vssd1 vccd1 vccd1 _16790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4089 _17719_/Q vssd1 vssd1 vccd1 vccd1 hold4089/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3344 _17678_/Q vssd1 vssd1 vccd1 vccd1 hold3344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2610 _14127_/X vssd1 vssd1 vccd1 vccd1 _17867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3355 _17080_/Q vssd1 vssd1 vccd1 vccd1 _11768_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3366 _17227_/Q vssd1 vssd1 vccd1 vccd1 hold3366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 _14019_/X vssd1 vssd1 vccd1 vccd1 _17815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ hold8/X _16106_/Q _08993_/S vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__mux2_1
Xhold2632 _14211_/X vssd1 vssd1 vccd1 vccd1 _17908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3377 _11578_/X vssd1 vssd1 vccd1 vccd1 _17016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkbuf_4
Xhold2643 _18308_/Q vssd1 vssd1 vccd1 vccd1 hold2643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3388 _16445_/Q vssd1 vssd1 vccd1 vccd1 hold3388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3399 _09682_/X vssd1 vssd1 vccd1 vccd1 _16384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2654 _15724_/Q vssd1 vssd1 vccd1 vccd1 hold2654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1920 _15607_/Q vssd1 vssd1 vccd1 vccd1 hold1920/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18458_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2665 _14293_/X vssd1 vssd1 vccd1 vccd1 _17946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 _08091_/X vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _15551_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07928_/X sky130_fd_sc_hd__or2_1
Xhold2676 _17861_/Q vssd1 vssd1 vccd1 vccd1 hold2676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__buf_4
Xhold1942 _14047_/X vssd1 vssd1 vccd1 vccd1 _17829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 _15573_/Q vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _14723_/X vssd1 vssd1 vccd1 vccd1 _18153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _09115_/X vssd1 vssd1 vccd1 vccd1 _16172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 _15567_/Q vssd1 vssd1 vccd1 vccd1 hold1964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1975 _16193_/Q vssd1 vssd1 vccd1 vccd1 hold1975/X sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _15537_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07859_/X sky130_fd_sc_hd__or2_1
Xhold1986 _15544_/X vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1997 _14787_/X vssd1 vssd1 vccd1 vccd1 _18184_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10870_ hold3985/X _11150_/B _10869_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10870_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09529_ hold3859/X _10001_/B _09528_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _09529_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _12933_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _17356_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ hold81/X _08598_/B _08999_/B _12470_/X _15414_/A vssd1 vssd1 vccd1 vccd1
+ hold82/A sky130_fd_sc_hd__o311a_1
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14210_ hold800/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__or2_1
X_11422_ hold3442/X _12320_/B _11421_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15190_ hold2943/X _15221_/B _15189_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ hold5949/X hold587/X _14140_/X _13925_/A vssd1 vssd1 vccd1 vccd1 hold588/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ hold4244/X _11735_/B _11352_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10304_ hold2306/X hold4706/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__mux2_1
X_14072_ _15199_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14072_/X sky130_fd_sc_hd__or2_1
X_11284_ hold5747/X _11789_/B _11283_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o211a_1
X_13023_ _17518_/Q hold901/X vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__or2_1
Xhold5280 _12340_/Y vssd1 vssd1 vccd1 vccd1 _17270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17900_ _17900_/CLK hold468/X vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_1
X_10235_ hold2115/X _16569_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__mux2_1
Xhold5291 _16340_/Q vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4590 _13393_/X vssd1 vssd1 vccd1 vccd1 _17584_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17831_ _17895_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_1
X_10166_ hold2592/X hold3699/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__mux2_1
X_17762_ _17890_/CLK _17762_/D vssd1 vssd1 vccd1 vccd1 _17762_/Q sky130_fd_sc_hd__dfxtp_1
X_10097_ hold2785/X hold3144/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__mux2_1
X_14974_ hold667/X _15018_/B vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__or2_1
X_16713_ _18047_/CLK _16713_/D vssd1 vssd1 vccd1 vccd1 _16713_/Q sky130_fd_sc_hd__dfxtp_1
X_13925_ _13925_/A hold438/X vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__and2_1
X_17693_ _17693_/CLK _17693_/D vssd1 vssd1 vccd1 vccd1 _17693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13856_ _17739_/Q _13856_/B _13865_/C vssd1 vssd1 vccd1 vccd1 _13856_/X sky130_fd_sc_hd__and3_1
X_16644_ _18204_/CLK _16644_/D vssd1 vssd1 vccd1 vccd1 _16644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _12813_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _17445_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _18131_/CLK _16575_/D vssd1 vssd1 vccd1 vccd1 _16575_/Q sky130_fd_sc_hd__dfxtp_1
X_13787_ hold1604/X hold5205/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13788_/B sky130_fd_sc_hd__mux2_1
X_10999_ hold4115/X _11216_/B _10998_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18314_ _18334_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 hold485/A sky130_fd_sc_hd__dfxtp_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12756_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _17422_/D sky130_fd_sc_hd__and2_1
X_15526_ hold2443/X _15560_/A2 _15525_/X _12885_/A vssd1 vssd1 vccd1 vccd1 _15526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15457_ hold400/X _09392_/C _09386_/D hold709/X _15456_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/B sky130_fd_sc_hd__a221o_1
X_18245_ _18422_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ _12885_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _17399_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14408_ hold2949/X hold209/X _14407_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18405_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15388_ hold531/X _09386_/A _09392_/D hold596/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18176_ _18176_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17127_ _17221_/CLK _17127_/D vssd1 vssd1 vccd1 vccd1 _17127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ hold2096/X _14326_/B _14338_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14339_/X
+ sky130_fd_sc_hd__o211a_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold516 hold516/A vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 hold527/A vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold538 hold538/A vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17058_ _17208_/CLK _17058_/D vssd1 vssd1 vccd1 vccd1 _17058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold549 hold549/A vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
X_16009_ _18416_/CLK _16009_/D vssd1 vssd1 vccd1 vccd1 _16009_/Q sky130_fd_sc_hd__dfxtp_1
X_08900_ hold179/X hold568/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__mux2_1
X_09880_ hold4753/X _10070_/B _09879_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09880_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08831_ _15304_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _16034_/D sky130_fd_sc_hd__and2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _14181_/X vssd1 vssd1 vccd1 vccd1 _17893_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _15568_/Q vssd1 vssd1 vccd1 vccd1 hold1216/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _15344_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__and2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _15750_/Q vssd1 vssd1 vccd1 vccd1 hold1227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _09083_/X vssd1 vssd1 vccd1 vccd1 _16156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _17870_/Q vssd1 vssd1 vccd1 vccd1 hold1249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08693_ hold71/X hold559/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09314_ hold1781/X _09325_/B _09313_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ _15521_/A hold2841/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09246_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09176_ _15559_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _13925_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08058_ _15517_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3130 _11172_/Y vssd1 vssd1 vccd1 vccd1 _11173_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10020_ _13166_/A _09924_/A _10019_/X vssd1 vssd1 vccd1 vccd1 _10020_/Y sky130_fd_sc_hd__a21oi_1
Xhold3141 _17100_/Q vssd1 vssd1 vccd1 vccd1 hold3141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3152 _13810_/Y vssd1 vssd1 vccd1 vccd1 _17723_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3163 _12366_/Y vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3174 _17108_/Q vssd1 vssd1 vccd1 vccd1 hold3174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3185 _17589_/Q vssd1 vssd1 vccd1 vccd1 hold3185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2440 _14965_/X vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2451 _16154_/Q vssd1 vssd1 vccd1 vccd1 hold2451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3196 _17576_/Q vssd1 vssd1 vccd1 vccd1 hold3196/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2462 _16181_/Q vssd1 vssd1 vccd1 vccd1 hold2462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2473 _18267_/Q vssd1 vssd1 vccd1 vccd1 hold2473/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 _09316_/X vssd1 vssd1 vccd1 vccd1 _16268_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2495 _15781_/Q vssd1 vssd1 vccd1 vccd1 hold2495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1750 _17898_/Q vssd1 vssd1 vccd1 vccd1 hold1750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 _15536_/X vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ hold4712/X _12311_/B _11970_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _11971_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1772 _07811_/X vssd1 vssd1 vccd1 vccd1 hold1772/X sky130_fd_sc_hd__buf_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _18079_/Q vssd1 vssd1 vccd1 vccd1 hold1783/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _13710_/A _13710_/B vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__or2_1
Xhold1794 _18076_/Q vssd1 vssd1 vccd1 vccd1 hold1794/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ hold2947/X hold3991/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__mux2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _15191_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__or2_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ _13737_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _13641_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ hold2729/X hold3892/X _11726_/C vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _18273_/CLK _16360_/D vssd1 vssd1 vccd1 vccd1 _16360_/Q sky130_fd_sc_hd__dfxtp_1
X_13572_ _13764_/A _13572_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ hold2601/X hold3974/X _11747_/C vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _16295_/Q _09362_/A _09392_/B hold532/X _15310_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/D sky130_fd_sc_hd__a221o_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ hold683/X hold3436/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__mux2_1
X_16291_ _18460_/CLK _16291_/D vssd1 vssd1 vccd1 vccd1 _16291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15242_ _15489_/A _15242_/B _15242_/C _15242_/D vssd1 vssd1 vccd1 vccd1 _15242_/X
+ sky130_fd_sc_hd__or4_1
X_18030_ _18054_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_28__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_28__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_12454_ _17320_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__or2_1
X_11405_ hold1357/X hold5677/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__mux2_1
X_15173_ hold770/X _15179_/B vssd1 vssd1 vccd1 vccd1 _15173_/X sky130_fd_sc_hd__or2_1
X_12385_ hold407/X _17286_/Q _12439_/S vssd1 vssd1 vccd1 vccd1 hold408/A sky130_fd_sc_hd__mux2_1
XFILLER_0_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ _14517_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14124_/X sky130_fd_sc_hd__or2_1
X_11336_ hold1679/X hold4619/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _14735_/A hold272/X vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__or2_4
X_11267_ hold2850/X hold3645/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__mux2_1
X_13006_ hold1089/X _13003_/Y _13005_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13006_/X
+ sky130_fd_sc_hd__o211a_1
X_10218_ _10524_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__or2_1
X_11198_ _16890_/Q _11213_/B _11213_/C vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_190_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18236_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17814_ _17877_/CLK _17814_/D vssd1 vssd1 vccd1 vccd1 _17814_/Q sky130_fd_sc_hd__dfxtp_1
X_10149_ _10515_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17745_ _17745_/CLK _17745_/D vssd1 vssd1 vccd1 vccd1 _17745_/Q sky130_fd_sc_hd__dfxtp_1
X_14957_ hold1580/X _14952_/B _14956_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _14957_/X
+ sky130_fd_sc_hd__o211a_1
X_13908_ _14517_/A hold1183/X hold244/X vssd1 vssd1 vccd1 vccd1 _13908_/X sky130_fd_sc_hd__mux2_1
X_17676_ _17708_/CLK _17676_/D vssd1 vssd1 vccd1 vccd1 _17676_/Q sky130_fd_sc_hd__dfxtp_1
X_14888_ _15227_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__or2_1
X_16627_ _18185_/CLK _16627_/D vssd1 vssd1 vccd1 vccd1 _16627_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ hold3846/X _13770_/A _13838_/X vssd1 vssd1 vccd1 vccd1 _13839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16558_ _18265_/CLK _16558_/D vssd1 vssd1 vccd1 vccd1 _16558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ hold944/X _15559_/B vssd1 vssd1 vccd1 vccd1 hold945/A sky130_fd_sc_hd__or2_1
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ _18243_/CLK _16489_/D vssd1 vssd1 vccd1 vccd1 _16489_/Q sky130_fd_sc_hd__dfxtp_1
X_09030_ hold179/X _16132_/Q _09056_/S vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__mux2_1
XFILLER_0_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18228_ _18228_/CLK hold856/X vssd1 vssd1 vccd1 vccd1 hold855/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18159_ _18183_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__buf_8
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold346 hold442/X vssd1 vssd1 vccd1 vccd1 hold443/A sky130_fd_sc_hd__clkbuf_2
Xhold357 hold28/X vssd1 vssd1 vccd1 vccd1 input25/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_278_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17889_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ hold1540/X _16468_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold379 input26/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__buf_1
XFILLER_0_159_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout804 _15066_/A vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_207_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17769_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout815 fanout816/X vssd1 vssd1 vccd1 vccd1 _14939_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout826 _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/C1 sky130_fd_sc_hd__buf_4
X_09863_ hold806/X hold3388/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__mux2_1
Xfanout837 _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14889_/C1 sky130_fd_sc_hd__clkbuf_8
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout848 _12331_/A vssd1 vssd1 vccd1 vccd1 _12343_/A sky130_fd_sc_hd__buf_6
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 hold5878/X vssd1 vssd1 vccd1 vccd1 _13312_/B1 sky130_fd_sc_hd__buf_6
X_08814_ hold41/X hold348/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__mux2_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _17960_/Q vssd1 vssd1 vccd1 vccd1 hold1002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 _13036_/X vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 _15823_/Q vssd1 vssd1 vccd1 vccd1 hold1024/X sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _18335_/Q _16422_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__mux2_1
Xhold1035 _17808_/Q vssd1 vssd1 vccd1 vccd1 hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1046 hold881/X vssd1 vssd1 vccd1 vccd1 input68/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ hold47/X _15993_/Q _08787_/S vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__mux2_1
Xhold1057 hold1298/X vssd1 vssd1 vccd1 vccd1 hold1057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _09288_/X vssd1 vssd1 vccd1 vccd1 _16254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _17834_/Q vssd1 vssd1 vccd1 vccd1 hold1079/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08676_ _09003_/A _08676_/B vssd1 vssd1 vccd1 vccd1 _15959_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _15557_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ hold2228/X _09164_/B _09158_/Y _14360_/A vssd1 vssd1 vccd1 vccd1 _09159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12170_ hold1134/X hold4671/X _13871_/C vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 hold880/A vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 hold891/A vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__buf_8
XFILLER_0_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11052_ _11061_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__or2_1
X_10003_ _11203_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10003_/Y sky130_fd_sc_hd__nor2_1
X_15860_ _17728_/CLK _15860_/D vssd1 vssd1 vccd1 vccd1 _15860_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2270 _17904_/Q vssd1 vssd1 vccd1 vccd1 hold2270/X sky130_fd_sc_hd__dlygate4sd3_1
X_14811_ hold2180/X _14822_/B _14810_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14811_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2281 _15850_/Q vssd1 vssd1 vccd1 vccd1 hold2281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2292 _07860_/X vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _17693_/CLK _15791_/D vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1580 _18265_/Q vssd1 vssd1 vccd1 vccd1 hold1580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17530_ _17530_/CLK _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _15189_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__or2_1
X_11954_ hold1958/X _17142_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__mux2_1
Xhold1591 hold6010/X vssd1 vssd1 vccd1 vccd1 _09456_/C sky130_fd_sc_hd__clkbuf_2
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _11103_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__or2_1
X_14673_ hold1905/X _14666_/B _14672_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14673_/X
+ sky130_fd_sc_hd__o211a_1
X_17461_ _18441_/CLK _17461_/D vssd1 vssd1 vccd1 vccd1 _17461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ hold1876/X hold3162/X _12368_/C vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16412_ _18389_/CLK _16412_/D vssd1 vssd1 vccd1 vccd1 _16412_/Q sky130_fd_sc_hd__dfxtp_1
X_13624_ hold4226/X _13814_/B _13623_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13624_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _11670_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17392_ _18454_/CLK _17392_/D vssd1 vssd1 vccd1 vccd1 _17392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16343_ _18360_/CLK _16343_/D vssd1 vssd1 vccd1 vccd1 _16343_/Q sky130_fd_sc_hd__dfxtp_1
X_13555_ hold4873/X _13859_/B _13554_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13555_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10767_ _11061_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12506_ _17346_/Q _12506_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16274_ _17375_/CLK _16274_/D vssd1 vssd1 vccd1 vccd1 _16274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ hold3552/X _13847_/B _13485_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _11082_/A _10698_/B vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _15225_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__or2_1
X_18013_ _18013_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
X_12437_ hold359/X hold387/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15156_ hold1763/X _15161_/B _15155_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _15156_/X
+ sky130_fd_sc_hd__o211a_1
X_12368_ _17280_/Q _12374_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and3_1
XFILLER_0_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14107_ hold2054/X _14094_/B _14106_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14107_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11319_ _12153_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__or2_1
X_15087_ _15195_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15087_/X sky130_fd_sc_hd__or2_1
X_12299_ _17257_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_300_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17730_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14038_ _15545_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15989_ _17343_/CLK _15989_/D vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__dfxtp_1
X_08530_ _13056_/C _17520_/Q _08868_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__or3_1
X_17728_ _17728_/CLK _17728_/D vssd1 vssd1 vccd1 vccd1 _17728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08461_ hold2435/X _08488_/B _08460_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17659_ _17691_/CLK _17659_/D vssd1 vssd1 vccd1 vccd1 _17659_/Q sky130_fd_sc_hd__dfxtp_1
X_08392_ hold624/A hold279/X hold298/A hold606/A vssd1 vssd1 vccd1 vccd1 _15508_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _09021_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _16123_/D sky130_fd_sc_hd__and2_1
XFILLER_0_170_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5802 hold5930/X vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5813 hold5813/A vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5824 _18410_/Q vssd1 vssd1 vccd1 vccd1 hold5824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold110 input28/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__buf_1
Xhold5835 hold5938/X vssd1 vssd1 vccd1 vccd1 hold5835/X sky130_fd_sc_hd__clkbuf_2
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__clkbuf_2
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5846 hold5939/X vssd1 vssd1 vccd1 vccd1 hold5846/X sky130_fd_sc_hd__clkbuf_2
Xhold5857 hold5857/A vssd1 vssd1 vccd1 vccd1 hold5857/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold143 hold172/X vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__buf_6
Xhold5868 _16284_/Q vssd1 vssd1 vccd1 vccd1 hold5868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5879 _07826_/X vssd1 vssd1 vccd1 vccd1 hold5879/X sky130_fd_sc_hd__buf_1
Xhold154 input22/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__buf_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 data_in[15] vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold187 hold248/X vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _12589_/S vssd1 vssd1 vccd1 vccd1 _12982_/S sky130_fd_sc_hd__clkbuf_8
Xfanout612 _09360_/Y vssd1 vssd1 vccd1 vccd1 _09362_/C sky130_fd_sc_hd__clkbuf_8
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09918_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__or2_1
Xfanout623 _09349_/Y vssd1 vssd1 vccd1 vccd1 _15485_/A2 sky130_fd_sc_hd__buf_6
Xfanout634 fanout660/X vssd1 vssd1 vccd1 vccd1 _12813_/A sky130_fd_sc_hd__clkbuf_4
Xfanout645 _12831_/A vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__buf_4
Xfanout656 fanout660/X vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__clkbuf_4
X_09846_ _09954_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__or2_1
XFILLER_0_176_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout667 fanout842/X vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout678 _14492_/C1 vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__buf_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _12951_/A vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__buf_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09951_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _09021_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _15985_/D sky130_fd_sc_hd__and2_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ hold14/X hold531/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__mux2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ _10651_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ hold2979/X hold3687/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13341_/B sky130_fd_sc_hd__mux2_1
X_10552_ hold4097/X _10589_/B _10551_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13311_/A1 _13269_/X _13270_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13271_/X
+ sky130_fd_sc_hd__o211a_2
X_10483_ hold4512/X _10073_/B _10482_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10483_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_129_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18389_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15010_ _15225_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _15010_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _12267_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12153_ _12153_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ hold5659/X _11213_/B _11103_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _11104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12084_ _12282_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__or2_1
X_16961_ _17873_/CLK _16961_/D vssd1 vssd1 vccd1 vccd1 _16961_/Q sky130_fd_sc_hd__dfxtp_1
X_15912_ _17287_/CLK _15912_/D vssd1 vssd1 vccd1 vccd1 hold719/A sky130_fd_sc_hd__dfxtp_1
X_11035_ hold5685/X _11765_/B _11034_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16892_ _18063_/CLK _16892_/D vssd1 vssd1 vccd1 vccd1 _16892_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _17734_/CLK _15843_/D vssd1 vssd1 vccd1 vccd1 _15843_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _17693_/CLK _15774_/D vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfxtp_1
X_12986_ hold3426/X _12985_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__mux2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17513_ _17513_/CLK _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14725_ hold1538/X _14718_/B _14724_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14725_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _12093_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__or2_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17444_ _17447_/CLK _17444_/D vssd1 vssd1 vccd1 vccd1 _17444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ _15103_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__or2_1
X_11868_ _12255_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13607_ _15789_/Q hold3212/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__mux2_1
X_10819_ hold4119/X _11177_/B _10818_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17375_ _17375_/CLK _17375_/D vssd1 vssd1 vccd1 vccd1 _17375_/Q sky130_fd_sc_hd__dfxtp_1
X_14587_ hold2872/X _14610_/B _14586_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ hold3841/X _12153_/A _11798_/X vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16326_ _18339_/CLK _16326_/D vssd1 vssd1 vccd1 vccd1 _16326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ _15818_/Q _17633_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13469_ hold2572/X hold5164/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13470_/B sky130_fd_sc_hd__mux2_1
X_16257_ _17487_/CLK _16257_/D vssd1 vssd1 vccd1 vccd1 _16257_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5109 _10909_/X vssd1 vssd1 vccd1 vccd1 _16793_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15208_ hold1401/X _15219_/B _15207_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _15208_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4408 _10117_/X vssd1 vssd1 vccd1 vccd1 _16529_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16188_ _18432_/CLK _16188_/D vssd1 vssd1 vccd1 vccd1 _16188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4419 _17006_/Q vssd1 vssd1 vccd1 vccd1 hold4419/X sky130_fd_sc_hd__dlygate4sd3_1
X_15139_ _15193_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15139_/X sky130_fd_sc_hd__or2_1
Xhold3707 _11221_/Y vssd1 vssd1 vccd1 vccd1 _16897_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3718 _10057_/Y vssd1 vssd1 vccd1 vccd1 _16509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3729 _10641_/Y vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07961_ hold1954/X _07991_/A2 _07960_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07961_/X
+ sky130_fd_sc_hd__o211a_1
X_09700_ hold5530/X _10780_/A2 _09699_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _09700_/X
+ sky130_fd_sc_hd__o211a_1
X_07892_ _14850_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__or2_1
X_09631_ hold3762/X _10028_/B _09630_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09631_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ hold5056/X _10571_/B _09561_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _09562_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08513_ _15517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__or2_1
X_09493_ _09494_/A _13055_/C _09494_/C vssd1 vssd1 vccd1 vccd1 _09493_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ hold1513/X _08433_/B _08443_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08375_ _09272_/A hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_293_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17252_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_222_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17907_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5610 _16464_/Q vssd1 vssd1 vccd1 vccd1 hold5610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5621 _16779_/Q vssd1 vssd1 vccd1 vccd1 hold5621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5632 _09928_/X vssd1 vssd1 vccd1 vccd1 _16466_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5643 _16432_/Q vssd1 vssd1 vccd1 vccd1 hold5643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5654 _11656_/X vssd1 vssd1 vccd1 vccd1 _17042_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4920 _11893_/X vssd1 vssd1 vccd1 vccd1 _17121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5665 _09889_/X vssd1 vssd1 vccd1 vccd1 _16453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5676 _16325_/Q vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4931 _17621_/Q vssd1 vssd1 vccd1 vccd1 hold4931/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4942 _11419_/X vssd1 vssd1 vccd1 vccd1 _16963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5687 _16794_/Q vssd1 vssd1 vccd1 vccd1 hold5687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4953 _17277_/Q vssd1 vssd1 vccd1 vccd1 hold4953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5698 _11380_/X vssd1 vssd1 vccd1 vccd1 _16950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4964 _11323_/X vssd1 vssd1 vccd1 vccd1 _16931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4975 _17608_/Q vssd1 vssd1 vccd1 vccd1 hold4975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4986 _12034_/X vssd1 vssd1 vccd1 vccd1 _17168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout420 _14054_/Y vssd1 vssd1 vccd1 vccd1 _14105_/A2 sky130_fd_sc_hd__buf_6
Xfanout431 _13173_/S vssd1 vssd1 vccd1 vccd1 _13309_/S sky130_fd_sc_hd__buf_8
Xhold4997 _17273_/Q vssd1 vssd1 vccd1 vccd1 hold4997/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout442 _13862_/C vssd1 vssd1 vccd1 vccd1 _13832_/C sky130_fd_sc_hd__buf_6
Xfanout453 _11741_/C vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__clkbuf_8
Xfanout464 fanout484/X vssd1 vssd1 vccd1 vccd1 _12332_/C sky130_fd_sc_hd__buf_4
Xfanout475 _11210_/C vssd1 vssd1 vccd1 vccd1 _11762_/C sky130_fd_sc_hd__clkbuf_8
Xfanout486 _10763_/S vssd1 vssd1 vccd1 vccd1 _11156_/C sky130_fd_sc_hd__clkbuf_8
X_09829_ hold5415/X _10025_/B _09828_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09829_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout497 fanout523/X vssd1 vssd1 vccd1 vccd1 _10763_/S sky130_fd_sc_hd__buf_4
X_12840_ _12843_/A _12840_/B vssd1 vssd1 vccd1 vccd1 _17456_/D sky130_fd_sc_hd__and2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12771_ _12804_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _17433_/D sky130_fd_sc_hd__and2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _12301_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11722_/Y sky130_fd_sc_hd__nor2_1
X_14510_ hold2866/X _14554_/A2 _14509_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14510_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15490_ _15490_/A1 _15483_/X _15489_/X _15490_/B1 hold5873/A vssd1 vssd1 vccd1 vccd1
+ _15490_/X sky130_fd_sc_hd__a32o_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ hold4075/X _11747_/B _11652_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11653_/X
+ sky130_fd_sc_hd__o211a_1
X_14441_ _14728_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14441_/X sky130_fd_sc_hd__or2_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _16692_/Q _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__and3_1
X_17160_ _17724_/CLK _17160_/D vssd1 vssd1 vccd1 vccd1 _17160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14372_ _15036_/A hold912/X vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ hold4113/X _12338_/B _11583_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16111_ _17341_/CLK _16111_/D vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__dfxtp_1
X_13323_ _13710_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ hold989/X hold4147/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__mux2_1
X_17091_ _17907_/CLK _17091_/D vssd1 vssd1 vccd1 vccd1 _17091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _18414_/CLK _16042_/D vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__dfxtp_1
X_13254_ _13254_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ hold1152/X _16646_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ hold4809/X _12299_/B _12204_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _12205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13185_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ hold2149/X hold4125/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__mux2_1
X_12136_ hold4502/X _13871_/B _12135_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12136_/X
+ sky130_fd_sc_hd__o211a_1
X_17993_ _18065_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
X_12067_ hold5023/X _12311_/B _12066_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o211a_1
X_16944_ _17855_/CLK _16944_/D vssd1 vssd1 vccd1 vccd1 _16944_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18416_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11018_ hold2717/X _16830_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11019_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17879_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16875_ _18046_/CLK _16875_/D vssd1 vssd1 vccd1 vccd1 _16875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _17649_/CLK _15826_/D vssd1 vssd1 vccd1 vccd1 _15826_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _17708_/CLK _15757_/D vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _14364_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _17499_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ _15209_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14708_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15688_ _17742_/CLK _15688_/D vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17427_ _17629_/CLK _17427_/D vssd1 vssd1 vccd1 vccd1 _17427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14639_ hold3105/X _14666_/B _14638_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08160_ hold892/X _15718_/Q _08170_/S vssd1 vssd1 vccd1 vccd1 hold893/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ _17487_/CLK _17358_/D vssd1 vssd1 vccd1 vccd1 _17358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16309_ _16314_/CLK _16309_/D vssd1 vssd1 vccd1 vccd1 _16309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ hold1930/X _08088_/B _08090_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17289_ _17289_/CLK _17289_/D vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4205 _17002_/Q vssd1 vssd1 vccd1 vccd1 hold4205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4216 _11665_/X vssd1 vssd1 vccd1 vccd1 _17045_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4227 _13624_/X vssd1 vssd1 vccd1 vccd1 _17661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4238 _17697_/Q vssd1 vssd1 vccd1 vccd1 hold4238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3504 _17626_/Q vssd1 vssd1 vccd1 vccd1 hold3504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4249 _10843_/X vssd1 vssd1 vccd1 vccd1 _16771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3515 _17268_/Q vssd1 vssd1 vccd1 vccd1 hold3515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3526 _17653_/Q vssd1 vssd1 vccd1 vccd1 hold3526/X sky130_fd_sc_hd__dlygate4sd3_1
X_08993_ hold380/X hold453/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__mux2_1
Xhold3537 _16972_/Q vssd1 vssd1 vccd1 vccd1 hold3537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3548 _16442_/Q vssd1 vssd1 vccd1 vccd1 hold3548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2803 _18135_/Q vssd1 vssd1 vccd1 vccd1 hold2803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 _15748_/Q vssd1 vssd1 vccd1 vccd1 hold2814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3559 _10288_/X vssd1 vssd1 vccd1 vccd1 _16586_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 _14187_/X vssd1 vssd1 vccd1 vccd1 _17896_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07944_ _15513_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2836 _15619_/Q vssd1 vssd1 vccd1 vccd1 hold2836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 _14743_/X vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2858 _16158_/Q vssd1 vssd1 vccd1 vccd1 hold2858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 _14707_/X vssd1 vssd1 vccd1 vccd1 _18145_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07875_ _14726_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ hold952/X hold5598/X _11066_/S vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ hold1181/X _13182_/A _10025_/C vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ hold681/X _09477_/C _09477_/A vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08427_ _15000_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ _15527_/A hold2182/X hold122/X vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _15513_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10554_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5440 _09637_/X vssd1 vssd1 vccd1 vccd1 _16369_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5451 _10717_/X vssd1 vssd1 vccd1 vccd1 _16729_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _10521_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__or2_1
Xhold5462 _16757_/Q vssd1 vssd1 vccd1 vccd1 hold5462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5473 _12139_/X vssd1 vssd1 vccd1 vccd1 _17203_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5484 _16830_/Q vssd1 vssd1 vccd1 vccd1 hold5484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5495 _11308_/X vssd1 vssd1 vccd1 vccd1 _16926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4750 _11266_/X vssd1 vssd1 vccd1 vccd1 _16912_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10182_ _10563_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4761 _17250_/Q vssd1 vssd1 vccd1 vccd1 hold4761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4772 _10702_/X vssd1 vssd1 vccd1 vccd1 _16724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4783 _17605_/Q vssd1 vssd1 vccd1 vccd1 hold4783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4794 _11953_/X vssd1 vssd1 vccd1 vccd1 _17141_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout250 _13713_/A vssd1 vssd1 vccd1 vccd1 _13800_/A sky130_fd_sc_hd__buf_4
X_14990_ _15205_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__or2_1
Xfanout261 fanout299/X vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__buf_2
Xfanout272 fanout299/X vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__clkbuf_4
Xfanout283 _12279_/A vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__clkbuf_4
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _17778_/D sky130_fd_sc_hd__and2_1
Xfanout294 fanout298/X vssd1 vssd1 vccd1 vccd1 _11697_/A sky130_fd_sc_hd__clkbuf_4
X_16660_ _18266_/CLK _16660_/D vssd1 vssd1 vccd1 vccd1 _16660_/Q sky130_fd_sc_hd__dfxtp_1
X_13872_ hold3945/X _13392_/A _13871_/X vssd1 vssd1 vccd1 vccd1 _13872_/Y sky130_fd_sc_hd__a21oi_1
X_15611_ _17227_/CLK _15611_/D vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ hold2018/X hold3054/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12823_/X sky130_fd_sc_hd__mux2_1
X_16591_ _18149_/CLK _16591_/D vssd1 vssd1 vccd1 vccd1 _16591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18330_ _18330_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ hold2357/X _15547_/B _15541_/Y _12666_/A vssd1 vssd1 vccd1 vccd1 _15542_/X
+ sky130_fd_sc_hd__o211a_1
X_12754_ hold1407/X _17429_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__mux2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18261_ _18315_/CLK hold866/X vssd1 vssd1 vccd1 vccd1 hold865/A sky130_fd_sc_hd__dfxtp_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ hold1977/X _17059_/Q _12341_/C vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15473_ _15473_/A _15473_/B vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__and2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ hold2695/X hold3056/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18215_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17212_ _17276_/CLK _17212_/D vssd1 vssd1 vccd1 vccd1 _17212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11636_ hold871/X hold4813/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__mux2_1
X_14424_ hold2338/X _14433_/B _14423_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _14424_/X
+ sky130_fd_sc_hd__o211a_1
X_18192_ _18192_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17143_ _17779_/CLK _17143_/D vssd1 vssd1 vccd1 vccd1 _17143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11567_ hold2676/X _17013_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__mux2_1
X_14355_ hold949/X hold1118/X hold275/X vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _10542_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__or2_1
X_13306_ _17589_/Q _17123_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__mux2_1
Xhold709 hold709/A vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17074_ _17890_/CLK _17074_/D vssd1 vssd1 vccd1 vccd1 _17074_/Q sky130_fd_sc_hd__dfxtp_1
X_14286_ _15508_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14286_/Y sky130_fd_sc_hd__nor2_2
X_11498_ hold2503/X _16990_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__mux2_1
X_16025_ _17524_/CLK _16025_/D vssd1 vssd1 vccd1 vccd1 hold673/A sky130_fd_sc_hd__dfxtp_1
X_13237_ _13236_/X hold3745/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ _10554_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ _13161_/X _13167_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17539_/D sky130_fd_sc_hd__o21a_1
X_12119_ hold1826/X hold4965/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__mux2_1
X_13099_ _13098_/X hold5896/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux2_1
X_17976_ _18042_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1409 _15202_/X vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16927_ _17829_/CLK _16927_/D vssd1 vssd1 vccd1 vccd1 _16927_/Q sky130_fd_sc_hd__dfxtp_1
X_16858_ _18034_/CLK _16858_/D vssd1 vssd1 vccd1 vccd1 _16858_/Q sky130_fd_sc_hd__dfxtp_1
X_15809_ _17724_/CLK _15809_/D vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16789_ _18158_/CLK _16789_/D vssd1 vssd1 vccd1 vccd1 _16789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ hold1311/X _09338_/A2 _09329_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ _15537_/A hold2087/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18459_ _18462_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08212_ hold2085/X _08213_/B _08211_/Y _08349_/A vssd1 vssd1 vccd1 vccd1 _08212_/X
+ sky130_fd_sc_hd__o211a_1
X_09192_ _15521_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08143_ _08143_/A hold197/X vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__and2_1
XFILLER_0_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08074_ _15533_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4002 _11392_/X vssd1 vssd1 vccd1 vccd1 _16954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4013 _10864_/X vssd1 vssd1 vccd1 vccd1 _16778_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4024 _17190_/Q vssd1 vssd1 vccd1 vccd1 hold4024/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4035 _16763_/Q vssd1 vssd1 vccd1 vccd1 hold4035/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3301 _17485_/Q vssd1 vssd1 vccd1 vccd1 hold3301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4046 _10774_/X vssd1 vssd1 vccd1 vccd1 _16748_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4057 _16661_/Q vssd1 vssd1 vccd1 vccd1 hold4057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3312 _10366_/X vssd1 vssd1 vccd1 vccd1 _16612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3323 _13576_/X vssd1 vssd1 vccd1 vccd1 _17645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4068 _13534_/X vssd1 vssd1 vccd1 vccd1 _17631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3334 _16589_/Q vssd1 vssd1 vccd1 vccd1 hold3334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4079 _16652_/Q vssd1 vssd1 vccd1 vccd1 hold4079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3345 _13579_/X vssd1 vssd1 vccd1 vccd1 _17646_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2600 _09151_/X vssd1 vssd1 vccd1 vccd1 _16188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2611 _15715_/Q vssd1 vssd1 vccd1 vccd1 hold2611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3356 _11674_/X vssd1 vssd1 vccd1 vccd1 _17048_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__buf_4
Xhold2622 _15596_/Q vssd1 vssd1 vccd1 vccd1 hold2622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3367 _12115_/X vssd1 vssd1 vccd1 vccd1 _17195_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _12430_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _16105_/D sky130_fd_sc_hd__and2_1
Xhold3378 _16404_/Q vssd1 vssd1 vccd1 vccd1 hold3378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 _18272_/Q vssd1 vssd1 vccd1 vccd1 hold2633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2644 _16256_/Q vssd1 vssd1 vccd1 vccd1 hold2644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3389 _09769_/X vssd1 vssd1 vccd1 vccd1 _16413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1910 _14619_/X vssd1 vssd1 vccd1 vccd1 _18103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__buf_4
Xhold2655 _08176_/X vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ hold1920/X _07924_/B _07926_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _07927_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1921 _07927_/X vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2666 _17864_/Q vssd1 vssd1 vccd1 vccd1 hold2666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2677 _14115_/X vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 _18237_/Q vssd1 vssd1 vccd1 vccd1 hold1932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 _07856_/X vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _15631_/Q vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _15623_/Q vssd1 vssd1 vccd1 vccd1 hold1954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 _17920_/Q vssd1 vssd1 vccd1 vccd1 hold2699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _07844_/X vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ hold1736/X _07869_/B _07857_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _07858_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1976 _09161_/X vssd1 vssd1 vccd1 vccd1 _16193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 _15770_/Q vssd1 vssd1 vccd1 vccd1 hold1987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1998 _17849_/Q vssd1 vssd1 vccd1 vccd1 hold1998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _18462_/Q vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__inv_2
XFILLER_0_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09948_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__or2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09463_/C _09463_/D _09458_/Y vssd1 vssd1 vccd1 vccd1 _16313_/D sky130_fd_sc_hd__o21a_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _17328_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__or2_1
Xclkbuf_5_27__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_27__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11421_ _11649_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14140_ hold466/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14140_/X sky130_fd_sc_hd__or2_1
X_11352_ _11640_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11352_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ hold4125/X _10640_/B _10302_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14071_ hold1082/X _14105_/A2 _14070_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11283_ _11694_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__or2_1
Xhold5270 _10026_/Y vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__dlygate4sd3_1
X_13022_ _09494_/A hold901/X _11203_/A vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__a21oi_2
Xhold5281 _16914_/Q vssd1 vssd1 vccd1 vccd1 hold5281/X sky130_fd_sc_hd__dlygate4sd3_1
X_10234_ hold4203/X _10643_/B _10233_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10234_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5292 _10029_/Y vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4580 _11482_/X vssd1 vssd1 vccd1 vccd1 _16984_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17830_ _17862_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4591 _16758_/Q vssd1 vssd1 vccd1 vccd1 hold4591/X sky130_fd_sc_hd__dlygate4sd3_1
X_10165_ hold4033/X _10643_/B _10164_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10165_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3890 _17017_/Q vssd1 vssd1 vccd1 vccd1 hold3890/X sky130_fd_sc_hd__dlygate4sd3_1
X_17761_ _17827_/CLK _17761_/D vssd1 vssd1 vccd1 vccd1 _17761_/Q sky130_fd_sc_hd__dfxtp_1
X_14973_ hold2633/X _15006_/B _14972_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _14973_/X
+ sky130_fd_sc_hd__o211a_1
X_10096_ hold5154/X _11177_/B _10095_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10096_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712_ _18043_/CLK _16712_/D vssd1 vssd1 vccd1 vccd1 _16712_/Q sky130_fd_sc_hd__dfxtp_1
X_13924_ hold466/A _17770_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 hold438/A sky130_fd_sc_hd__mux2_1
X_17692_ _17692_/CLK _17692_/D vssd1 vssd1 vccd1 vccd1 _17692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16643_ _18230_/CLK _16643_/D vssd1 vssd1 vccd1 vccd1 _16643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _13888_/A _13855_/B vssd1 vssd1 vccd1 vccd1 _13855_/Y sky130_fd_sc_hd__nor2_1
X_12806_ hold3493/X _12805_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__mux2_1
X_16574_ _18222_/CLK _16574_/D vssd1 vssd1 vccd1 vccd1 _16574_/Q sky130_fd_sc_hd__dfxtp_1
X_13786_ hold5211/X _13883_/B _13785_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13786_/X
+ sky130_fd_sc_hd__o211a_1
X_10998_ _10998_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _10998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _18391_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _15525_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15525_/X sky130_fd_sc_hd__or2_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ hold3077/X _12736_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12738_/B sky130_fd_sc_hd__mux2_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18380_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
X_15456_ hold401/X _09365_/B _15487_/B1 _16098_/Q vssd1 vssd1 vccd1 vccd1 _15456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ hold3022/X _12667_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14407_ _14980_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18175_ _18267_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _12204_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15387_ hold445/X _15479_/A2 _09386_/D hold519/X _15386_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12599_ hold3216/X _12598_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17126_ _17592_/CLK _17126_/D vssd1 vssd1 vccd1 vccd1 _17126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14338_ _14786_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__or2_1
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold528 hold528/A vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold539 hold539/A vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _17777_/CLK _17057_/D vssd1 vssd1 vccd1 vccd1 _17057_/Q sky130_fd_sc_hd__dfxtp_1
X_14269_ hold2046/X _14272_/B _14268_/Y _14402_/C1 vssd1 vssd1 vccd1 vccd1 _14269_/X
+ sky130_fd_sc_hd__o211a_1
X_16008_ _18422_/CLK _16008_/D vssd1 vssd1 vccd1 vccd1 _16008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18241_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ hold59/X hold680/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__mux2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _15614_/Q vssd1 vssd1 vccd1 vccd1 hold1206/X sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ hold179/X hold308/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__mux2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _07846_/X vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _08231_/X vssd1 vssd1 vccd1 vccd1 _15750_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ _18055_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1239 _17763_/Q vssd1 vssd1 vccd1 vccd1 hold1239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08692_ _15304_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _15967_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _15535_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _12777_/A _09244_/B vssd1 vssd1 vccd1 vccd1 _16233_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ hold2767/X _09177_/A2 _09174_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08126_ _14866_/A hold1203/X hold196/X vssd1 vssd1 vccd1 vccd1 _08127_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08057_ hold1677/X _08082_/B _08056_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _08057_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3120 _17368_/Q vssd1 vssd1 vccd1 vccd1 hold3120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3131 _11173_/Y vssd1 vssd1 vccd1 vccd1 _16881_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3142 _12309_/Y vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3153 _17114_/Q vssd1 vssd1 vccd1 vccd1 hold3153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3164 _12367_/Y vssd1 vssd1 vccd1 vccd1 _17279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3175 _12333_/Y vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2430 _14281_/X vssd1 vssd1 vccd1 vccd1 _17941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3186 _13887_/Y vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2441 _15662_/Q vssd1 vssd1 vccd1 vccd1 hold2441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3197 _13848_/Y vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2452 _09079_/X vssd1 vssd1 vccd1 vccd1 _16154_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08959_ hold81/X hold725/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__mux2_1
Xhold2463 _09137_/X vssd1 vssd1 vccd1 vccd1 _16181_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 _14961_/X vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1740 _15678_/Q vssd1 vssd1 vccd1 vccd1 hold1740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 _17928_/Q vssd1 vssd1 vccd1 vccd1 hold2485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2496 _08296_/X vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1751 _14191_/X vssd1 vssd1 vccd1 vccd1 _17898_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _12267_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__or2_1
Xhold1762 _18432_/Q vssd1 vssd1 vccd1 vccd1 hold1762/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1773 _07812_/Y vssd1 vssd1 vccd1 vccd1 hold1773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _14568_/X vssd1 vssd1 vccd1 vccd1 hold1784/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10921_ hold4405/X _11222_/B _10920_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10921_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1795 _14562_/X vssd1 vssd1 vccd1 vccd1 hold1795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ hold2553/X hold4259/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ hold4921/X _10852_/A2 _10851_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ hold1387/X _17644_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ hold5679/X _11201_/B _10782_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ hold569/X _09367_/A _15446_/B1 hold567/X vssd1 vssd1 vccd1 vccd1 _15310_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _13002_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _17350_/D sky130_fd_sc_hd__and2_1
X_16290_ _16314_/CLK _16290_/D vssd1 vssd1 vccd1 vccd1 _16290_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15241_ _09404_/B _15477_/A2 _15487_/B1 hold458/X _15240_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/D sky130_fd_sc_hd__a221o_1
X_12453_ hold35/X _12509_/A2 _12505_/A3 _12452_/X _12422_/A vssd1 vssd1 vccd1 vccd1
+ hold36/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11404_ hold5486/X _12329_/B _11403_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12384_ _12430_/A _12384_/B vssd1 vssd1 vccd1 vccd1 _17285_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15172_ hold5982/X hold609/X _15171_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 hold610/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ hold2551/X hold587/X _14122_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14123_/X
+ sky130_fd_sc_hd__o211a_1
X_11335_ hold4947/X _12299_/B _11334_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11335_/X
+ sky130_fd_sc_hd__o211a_1
X_11266_ hold4749/X _12320_/B _11265_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o211a_1
X_14054_ _14735_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__nor2_1
X_10217_ hold2453/X _16563_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__mux2_1
X_13005_ _15183_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__or2_1
X_11197_ _12331_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/Y sky130_fd_sc_hd__nor2_1
X_17813_ _17877_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_1
X_10148_ hold2252/X _16540_/Q _10610_/C vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _17744_/CLK _17744_/D vssd1 vssd1 vccd1 vccd1 _17744_/Q sky130_fd_sc_hd__dfxtp_1
X_14956_ _15225_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__or2_1
X_10079_ _18075_/Q hold3431/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _14380_/A _13907_/B vssd1 vssd1 vccd1 vccd1 _17761_/D sky130_fd_sc_hd__and2_1
X_17675_ _17701_/CLK _17675_/D vssd1 vssd1 vccd1 vccd1 _17675_/Q sky130_fd_sc_hd__dfxtp_1
X_14887_ hold1582/X _14882_/B _14886_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16626_ _18216_/CLK _16626_/D vssd1 vssd1 vccd1 vccd1 _16626_/Q sky130_fd_sc_hd__dfxtp_1
X_13838_ _17733_/Q _13868_/B _13865_/C vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__and3_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ _18215_/CLK _16557_/D vssd1 vssd1 vccd1 vccd1 _16557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ hold1218/X hold3416/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15508_ _15508_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _15551_/B sky130_fd_sc_hd__or2_2
XFILLER_0_85_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16488_ _18273_/CLK _16488_/D vssd1 vssd1 vccd1 vccd1 _16488_/Q sky130_fd_sc_hd__dfxtp_1
X_18227_ _18227_/CLK hold990/X vssd1 vssd1 vccd1 vccd1 hold989/A sky130_fd_sc_hd__dfxtp_1
X_15439_ _15957_/Q _09386_/A _15437_/X vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18158_ _18158_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 hold25/X vssd1 vssd1 vccd1 vccd1 input33/A sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ _17779_/CLK _17109_/D vssd1 vssd1 vccd1 vccd1 _17109_/Q sky130_fd_sc_hd__dfxtp_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ _18217_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
Xhold336 hold336/A vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold358 input25/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ hold5514/X _10001_/B _09930_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold369 hold369/A vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout805 fanout816/X vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout816 fanout841/X vssd1 vssd1 vccd1 vccd1 fanout816/X sky130_fd_sc_hd__buf_4
X_09862_ hold5427/X _10013_/B _09861_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09862_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout827 _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14885_/C1 sky130_fd_sc_hd__buf_4
Xfanout838 _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/C1 sky130_fd_sc_hd__buf_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _11791_/A vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__buf_6
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _15454_/A _08813_/B vssd1 vssd1 vccd1 vccd1 _16025_/D sky130_fd_sc_hd__and2_1
Xhold1003 _14321_/X vssd1 vssd1 vccd1 vccd1 _17960_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ hold5352/X _10016_/B _09792_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09793_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _18440_/Q vssd1 vssd1 vccd1 vccd1 hold1014/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_247_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _15698_/Q vssd1 vssd1 vccd1 vccd1 hold1025/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _14005_/X vssd1 vssd1 vccd1 vccd1 _17808_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 input68/X vssd1 vssd1 vccd1 vccd1 hold882/A sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _12422_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _15992_/D sky130_fd_sc_hd__and2_1
Xhold1058 hold1058/A vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__buf_8
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 la_data_in[24] vssd1 vssd1 vccd1 vccd1 hold1069/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ hold41/X hold451/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08676_/B sky130_fd_sc_hd__mux2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ hold2652/X _09216_/B _09226_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09227_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ _15541_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09089_ hold2635/X _09119_/A2 _09088_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ hold2312/X _16864_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold870 hold870/A vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 hold881/A vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 hold892/A vssd1 vssd1 vccd1 vccd1 hold892/X sky130_fd_sc_hd__buf_8
X_11051_ hold954/X _16841_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__mux2_1
X_10002_ _13118_/A _09948_/A _10001_/X vssd1 vssd1 vccd1 vccd1 _10002_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2260 _15595_/Q vssd1 vssd1 vccd1 vccd1 hold2260/X sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ _14988_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__or2_1
Xhold2271 _14203_/X vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2282 _08440_/X vssd1 vssd1 vccd1 vccd1 _15850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2293 _18157_/Q vssd1 vssd1 vccd1 vccd1 hold2293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _17693_/CLK _15790_/D vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1570 _14458_/X vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 _14957_/X vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ hold2797/X _14774_/B _14740_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14741_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ hold4793/X _11798_/B _11952_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11953_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1592 _09413_/X vssd1 vssd1 vccd1 vccd1 _16292_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _18441_/CLK _17460_/D vssd1 vssd1 vccd1 vccd1 _17460_/Q sky130_fd_sc_hd__dfxtp_1
X_10904_ hold1989/X _16792_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10905_/B sky130_fd_sc_hd__mux2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14672_ _14726_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__or2_1
X_11884_ hold4423/X _13871_/B _11883_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o211a_1
X_16411_ _18396_/CLK _16411_/D vssd1 vssd1 vccd1 vccd1 _16411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13623_ _13800_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__or2_1
X_17391_ _18454_/CLK _17391_/D vssd1 vssd1 vccd1 vccd1 _17391_/Q sky130_fd_sc_hd__dfxtp_1
X_10835_ hold2596/X hold4211/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16342_ _18319_/CLK _16342_/D vssd1 vssd1 vccd1 vccd1 _16342_/Q sky130_fd_sc_hd__dfxtp_1
X_13554_ _13764_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__or2_1
X_10766_ hold1061/X _16746_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ hold62/X _12509_/A2 _12505_/A3 _12504_/X _12422_/A vssd1 vssd1 vccd1 vccd1
+ hold63/A sky130_fd_sc_hd__o311a_1
XFILLER_0_192_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16273_ _17375_/CLK _16273_/D vssd1 vssd1 vccd1 vccd1 _16273_/Q sky130_fd_sc_hd__dfxtp_1
X_13485_ _13758_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__or2_1
X_10697_ hold2940/X hold3648/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18012_ _18013_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ hold978/X _15219_/B _15223_/X _15026_/A vssd1 vssd1 vccd1 vccd1 hold979/A
+ sky130_fd_sc_hd__o211a_1
X_12436_ _15284_/A _12436_/B vssd1 vssd1 vccd1 vccd1 _17311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15155_ _15209_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12367_ _13888_/A _12367_/B vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ _14786_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__or2_1
X_11318_ hold2515/X hold3841/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__mux2_1
X_12298_ _13822_/A _12298_/B vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__nor2_1
X_15086_ hold2926/X _15109_/B _15085_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _15086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ hold1799/X _14036_/B _14036_/Y _14171_/C1 vssd1 vssd1 vccd1 vccd1 _14037_/X
+ sky130_fd_sc_hd__o211a_1
X_11249_ hold2874/X hold3737/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15988_ _17531_/CLK _15988_/D vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__dfxtp_1
X_17727_ _17730_/CLK _17727_/D vssd1 vssd1 vccd1 vccd1 _17727_/Q sky130_fd_sc_hd__dfxtp_1
X_14939_ hold1659/X _14946_/B _14938_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ _15519_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08460_/X sky130_fd_sc_hd__or2_1
X_17658_ _17693_/CLK _17658_/D vssd1 vssd1 vccd1 vccd1 _17658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _18231_/CLK _16609_/D vssd1 vssd1 vccd1 vccd1 _16609_/Q sky130_fd_sc_hd__dfxtp_1
X_08391_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _15827_/D sky130_fd_sc_hd__and2_1
X_17589_ _17749_/CLK _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ hold26/X hold374/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5803 output93/X vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_12
Xhold100 hold7/X vssd1 vssd1 vccd1 vccd1 input18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5814 hold6041/X vssd1 vssd1 vccd1 vccd1 hold5814/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5825 hold5825/A vssd1 vssd1 vccd1 vccd1 hold5825/X sky130_fd_sc_hd__buf_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5836 hold5836/A vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_12
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__clkbuf_16
Xhold5847 hold5847/A vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_12
Xhold133 data_in[11] vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5858 hold5942/X vssd1 vssd1 vccd1 vccd1 hold5858/X sky130_fd_sc_hd__buf_2
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5869 hold5869/A vssd1 vssd1 vccd1 vccd1 hold5869/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold177 hold10/X vssd1 vssd1 vccd1 vccd1 input11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold250/X vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__buf_2
XFILLER_0_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ hold1363/X hold3711/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__mux2_1
Xfanout602 hold2212/X vssd1 vssd1 vccd1 vccd1 _12679_/S sky130_fd_sc_hd__buf_4
Xfanout613 _09360_/Y vssd1 vssd1 vccd1 vccd1 _15486_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_186_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout624 _15484_/A2 vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__clkbuf_8
Xfanout635 _12777_/A vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout646 fanout660/X vssd1 vssd1 vccd1 vccd1 _12831_/A sky130_fd_sc_hd__buf_4
X_09845_ hold1714/X hold4607/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout657 _14360_/A vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__buf_4
Xfanout668 _08137_/A vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__buf_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout679 _14492_/C1 vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__buf_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ hold1684/X hold3398/X _10067_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__mux2_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ hold291/X hold389/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__mux2_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _12426_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _15951_/D sky130_fd_sc_hd__and2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _13002_/A _08589_/B vssd1 vssd1 vccd1 vccd1 _15918_/D sky130_fd_sc_hd__and2_1
XFILLER_0_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ hold3754/X _10422_/A _10619_/X vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ _10551_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _10506_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__or2_1
X_13270_ _13270_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ hold2256/X hold4785/X _12356_/C vssd1 vssd1 vccd1 vccd1 _12222_/B sky130_fd_sc_hd__mux2_1
X_12152_ hold2650/X hold4820/X _12152_/S vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_169_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18210_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11103_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12083_ hold2764/X hold4710/X _12377_/C vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__mux2_1
X_16960_ _17893_/CLK _16960_/D vssd1 vssd1 vccd1 vccd1 _16960_/Q sky130_fd_sc_hd__dfxtp_1
X_15911_ _18409_/CLK _15911_/D vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__dfxtp_1
X_11034_ _11670_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__or2_1
X_16891_ _18062_/CLK _16891_/D vssd1 vssd1 vccd1 vccd1 _16891_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _17701_/CLK hold834/X vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__dfxtp_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _18319_/Q vssd1 vssd1 vccd1 vccd1 hold2090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _17692_/CLK _15773_/D vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfxtp_1
X_12985_ hold2544/X hold3418/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__mux2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17512_ _17513_/CLK _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_1
X_14724_ _15225_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__or2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ hold1049/X hold4727/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__mux2_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17448_/CLK _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ hold1708/X _14666_/B _14654_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14655_/X
+ sky130_fd_sc_hd__o211a_1
X_11867_ hold2084/X hold3868/X _13388_/S vssd1 vssd1 vccd1 vccd1 _11868_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ hold4520/X _13814_/B _13605_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__o211a_1
X_17374_ _17375_/CLK _17374_/D vssd1 vssd1 vccd1 vccd1 _17374_/Q sky130_fd_sc_hd__dfxtp_1
X_10818_ _11082_/A _10818_/B vssd1 vssd1 vccd1 vccd1 _10818_/X sky130_fd_sc_hd__or2_1
X_14586_ _14980_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11798_ _17090_/Q _11798_/B _12152_/S vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__and3_1
X_16325_ _18304_/CLK _16325_/D vssd1 vssd1 vccd1 vccd1 _16325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13537_ hold4230/X _13832_/B _13536_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _11640_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ _17487_/CLK _16256_/D vssd1 vssd1 vccd1 vccd1 _16256_/Q sky130_fd_sc_hd__dfxtp_1
X_13468_ hold3550/X _13886_/B _13467_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15207_ _15207_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__or2_1
X_12419_ hold17/X hold326/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12420_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16187_ _18451_/CLK _16187_/D vssd1 vssd1 vccd1 vccd1 _16187_/Q sky130_fd_sc_hd__dfxtp_1
X_13399_ hold5082/X _13880_/B _13398_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13399_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4409 _17088_/Q vssd1 vssd1 vccd1 vccd1 hold4409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ hold1714/X hold609/X _15137_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15138_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3708 _16728_/Q vssd1 vssd1 vccd1 vccd1 hold3708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3719 _16906_/Q vssd1 vssd1 vccd1 vccd1 hold3719/X sky130_fd_sc_hd__dlygate4sd3_1
X_15069_ _15123_/A hold1277/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15070_/B sky130_fd_sc_hd__mux2_1
X_07960_ _15529_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07960_/X sky130_fd_sc_hd__or2_1
X_07891_ hold2870/X _07918_/B _07890_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07891_/X
+ sky130_fd_sc_hd__o211a_1
X_09630_ _09918_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _10380_/A _09561_/B vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__or2_1
X_08512_ hold1642/X _08503_/Y _08511_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _08512_/X
+ sky130_fd_sc_hd__o211a_1
X_09492_ _13030_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _09494_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ _15123_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08374_ hold86/X _15819_/Q hold122/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__mux2_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5600 _16457_/Q vssd1 vssd1 vccd1 vccd1 hold5600/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5611 _09826_/X vssd1 vssd1 vccd1 vccd1 _16432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5622 _10771_/X vssd1 vssd1 vccd1 vccd1 _16747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5633 _16946_/Q vssd1 vssd1 vccd1 vccd1 hold5633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5644 _09730_/X vssd1 vssd1 vccd1 vccd1 _16400_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4910 _12226_/X vssd1 vssd1 vccd1 vccd1 _17232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5655 _16356_/Q vssd1 vssd1 vccd1 vccd1 hold5655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5666 _16402_/Q vssd1 vssd1 vccd1 vccd1 hold5666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4921 _16806_/Q vssd1 vssd1 vccd1 vccd1 hold4921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4932 _13408_/X vssd1 vssd1 vccd1 vccd1 _17589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5677 _16959_/Q vssd1 vssd1 vccd1 vccd1 hold5677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4943 _17738_/Q vssd1 vssd1 vccd1 vccd1 hold4943/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_262_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5688 _10816_/X vssd1 vssd1 vccd1 vccd1 _16762_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4954 _12265_/X vssd1 vssd1 vccd1 vccd1 _17245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5699 _16368_/Q vssd1 vssd1 vccd1 vccd1 hold5699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4965 _17197_/Q vssd1 vssd1 vccd1 vccd1 hold4965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4976 _13369_/X vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout410 _14266_/B vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__buf_6
Xhold4987 _16710_/Q vssd1 vssd1 vccd1 vccd1 hold4987/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout421 _14050_/B vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout432 _13197_/S vssd1 vssd1 vccd1 vccd1 _13173_/S sky130_fd_sc_hd__buf_8
Xhold4998 _12253_/X vssd1 vssd1 vccd1 vccd1 _17241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout443 fanout484/X vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__clkbuf_8
Xfanout454 fanout484/X vssd1 vssd1 vccd1 vccd1 _11741_/C sky130_fd_sc_hd__buf_4
Xfanout465 _13886_/C vssd1 vssd1 vccd1 vccd1 _13883_/C sky130_fd_sc_hd__clkbuf_8
Xfanout476 _11672_/S vssd1 vssd1 vccd1 vccd1 _11210_/C sky130_fd_sc_hd__buf_4
X_09828_ _09924_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__or2_1
Xfanout487 _10874_/S vssd1 vssd1 vccd1 vccd1 _11066_/S sky130_fd_sc_hd__clkbuf_8
Xfanout498 _10562_/S vssd1 vssd1 vccd1 vccd1 _11177_/C sky130_fd_sc_hd__clkbuf_8
X_09759_ _09975_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__or2_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ hold3406/X _12769_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__mux2_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ hold3778/X _12204_/A _11720_/X vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ hold5979/X _14433_/B hold771/X _14376_/A vssd1 vssd1 vccd1 vccd1 hold772/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__or2_1
X_10603_ _10651_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10603_/Y sky130_fd_sc_hd__nor2_1
X_14371_ _15105_/A hold911/X hold275/X vssd1 vssd1 vccd1 vccd1 hold912/A sky130_fd_sc_hd__mux2_1
XFILLER_0_52_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _12051_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16110_ _17313_/CLK _16110_/D vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ hold1642/X hold3907/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__mux2_1
X_10534_ hold4581/X _10628_/B _10533_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10534_/X
+ sky130_fd_sc_hd__o211a_1
X_17090_ _17905_/CLK _17090_/D vssd1 vssd1 vccd1 vccd1 _17090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _18425_/CLK _16041_/D vssd1 vssd1 vccd1 vccd1 hold470/A sky130_fd_sc_hd__dfxtp_1
X_13253_ _13252_/X hold4003/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__mux2_1
X_10465_ hold3543/X _10465_/A2 _10464_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13184_ _13177_/X _13183_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17541_/D sky130_fd_sc_hd__o21a_1
X_10396_ hold3204/X _10649_/B _10395_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _13392_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__or2_1
X_17992_ _18158_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16943_ _17887_/CLK _16943_/D vssd1 vssd1 vccd1 vccd1 _16943_/Q sky130_fd_sc_hd__dfxtp_1
X_12066_ _13794_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ hold4475/X _11789_/B _11016_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16874_ _17981_/CLK _16874_/D vssd1 vssd1 vccd1 vccd1 _16874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15825_ _17738_/CLK _15825_/D vssd1 vssd1 vccd1 vccd1 _15825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _17701_/CLK _15756_/D vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12968_ hold3059/X _12967_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_66_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ hold2868/X _14718_/B _14706_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14707_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _13716_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__or2_1
X_15687_ _17211_/CLK _15687_/D vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ hold3121/X _12898_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17426_ _17629_/CLK _17426_/D vssd1 vssd1 vccd1 vccd1 _17426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ _15193_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17357_ _17487_/CLK _17357_/D vssd1 vssd1 vccd1 vccd1 _17357_/Q sky130_fd_sc_hd__dfxtp_1
X_14569_ _15193_/A _14557_/Y hold1784/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _16314_/CLK _16308_/D vssd1 vssd1 vccd1 vccd1 _16308_/Q sky130_fd_sc_hd__dfxtp_1
X_08090_ _15549_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08090_/X sky130_fd_sc_hd__or2_1
X_17288_ _17292_/CLK _17288_/D vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16239_ _17432_/CLK _16239_/D vssd1 vssd1 vccd1 vccd1 _16239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4206 _11440_/X vssd1 vssd1 vccd1 vccd1 _16970_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4217 _17253_/Q vssd1 vssd1 vccd1 vccd1 hold4217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4228 _16850_/Q vssd1 vssd1 vccd1 vccd1 hold4228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4239 _13636_/X vssd1 vssd1 vccd1 vccd1 _17665_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3505 _13423_/X vssd1 vssd1 vccd1 vccd1 _17594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3516 _12238_/X vssd1 vssd1 vccd1 vccd1 _17236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3527 _13504_/X vssd1 vssd1 vccd1 vccd1 _17621_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08992_ _12428_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _16113_/D sky130_fd_sc_hd__and2_1
Xhold3538 _11350_/X vssd1 vssd1 vccd1 vccd1 _16940_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3549 _09760_/X vssd1 vssd1 vccd1 vccd1 _16410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2804 _14687_/X vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 _08224_/X vssd1 vssd1 vccd1 vccd1 _15748_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07943_ hold1206/X _07991_/A2 _07942_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07943_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2826 _16155_/Q vssd1 vssd1 vccd1 vccd1 hold2826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2837 _07953_/X vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2848 _18059_/Q vssd1 vssd1 vccd1 vccd1 hold2848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2859 _09087_/X vssd1 vssd1 vccd1 vccd1 _16158_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07874_ hold1422/X _07869_/B _07873_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _07874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09613_ hold5516/X _09998_/B _09612_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09613_/X
+ sky130_fd_sc_hd__o211a_1
X_09544_ hold5639/X _10016_/B _09543_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ hold681/X _09477_/C _09474_/Y vssd1 vssd1 vccd1 vccd1 _16319_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_175_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ hold1114/X _08433_/B _08425_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_26__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_26__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ _08359_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _15810_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ hold1387/X _08336_/A2 _08287_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5430 _09913_/X vssd1 vssd1 vccd1 vccd1 _16461_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5441 _16882_/Q vssd1 vssd1 vccd1 vccd1 hold5441/X sky130_fd_sc_hd__dlygate4sd3_1
X_10250_ hold2157/X hold4273/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__mux2_1
Xhold5452 _16767_/Q vssd1 vssd1 vccd1 vccd1 hold5452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5463 _10705_/X vssd1 vssd1 vccd1 vccd1 _16725_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5474 _16895_/Q vssd1 vssd1 vccd1 vccd1 hold5474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4740 _12010_/X vssd1 vssd1 vccd1 vccd1 _17160_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5485 _10924_/X vssd1 vssd1 vccd1 vccd1 _16798_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10181_ hold2905/X _16551_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__mux2_1
Xhold4751 _16802_/Q vssd1 vssd1 vccd1 vccd1 hold4751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5496 _16456_/Q vssd1 vssd1 vccd1 vccd1 hold5496/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4762 _12184_/X vssd1 vssd1 vccd1 vccd1 _17218_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4773 _17278_/Q vssd1 vssd1 vccd1 vccd1 hold4773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4784 _13360_/X vssd1 vssd1 vccd1 vccd1 _17573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4795 _17143_/Q vssd1 vssd1 vccd1 vccd1 hold4795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout240 _09952_/A2 vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__clkbuf_4
Xfanout251 fanout299/X vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__clkbuf_4
Xfanout262 _11616_/A vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__clkbuf_4
Xfanout273 _13770_/A vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__buf_4
X_13940_ _14728_/A hold2515/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__mux2_1
Xfanout284 _12279_/A vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__buf_4
Xfanout295 _11031_/A vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__buf_4
X_13871_ _17744_/Q _13871_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _13871_/X sky130_fd_sc_hd__and3_1
X_15610_ _18445_/CLK _15610_/D vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfxtp_1
X_12822_ _12825_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _17450_/D sky130_fd_sc_hd__and2_1
XFILLER_0_186_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16590_ _18265_/CLK _16590_/D vssd1 vssd1 vccd1 vccd1 _16590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12753_ _12753_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _17427_/D sky130_fd_sc_hd__and2_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18396_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11704_ hold4583/X _11798_/B _11703_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11704_/X
+ sky130_fd_sc_hd__o211a_1
X_15472_ _15481_/A1 _15465_/X _15471_/X _15481_/B1 hold5871/A vssd1 vssd1 vccd1 vccd1
+ _15472_/X sky130_fd_sc_hd__a32o_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12684_ _12825_/A _12684_/B vssd1 vssd1 vccd1 vccd1 _17404_/D sky130_fd_sc_hd__and2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17211_/CLK _17211_/D vssd1 vssd1 vccd1 vccd1 _17211_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _15103_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14423_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18191_ _18223_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
X_11635_ hold4401/X _11732_/B _11634_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11635_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17142_ _17769_/CLK _17142_/D vssd1 vssd1 vccd1 vccd1 _17142_/Q sky130_fd_sc_hd__dfxtp_1
X_14354_ _14368_/A _14354_/B vssd1 vssd1 vccd1 vccd1 _17976_/D sky130_fd_sc_hd__and2_1
X_11566_ hold5367/X _11762_/B _11565_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_184_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18140_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13305_ _13305_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13305_/X sky130_fd_sc_hd__and2_1
X_10517_ hold2283/X hold3234/X _10523_/S vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17073_ _17889_/CLK _17073_/D vssd1 vssd1 vccd1 vccd1 _17073_/Q sky130_fd_sc_hd__dfxtp_1
X_14285_ hold5956/X _14266_/B hold785/X _14352_/A vssd1 vssd1 vccd1 vccd1 hold786/A
+ sky130_fd_sc_hd__o211a_1
X_11497_ hold5334/X _12329_/B _11496_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11497_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18371_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16024_ _17323_/CLK _16024_/D vssd1 vssd1 vccd1 vccd1 hold471/A sky130_fd_sc_hd__dfxtp_1
X_13236_ hold5297/X _13235_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10448_ hold1629/X _16640_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ _13183_/A1 _13165_/X _13166_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13167_/X
+ sky130_fd_sc_hd__o211a_1
X_10379_ hold2379/X hold3453/X _10568_/C vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12118_ hold4684/X _12308_/B _12117_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__o211a_1
X_13098_ _17563_/Q _17097_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
X_17975_ _18071_/CLK hold828/X vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ hold4653/X _12377_/B _12048_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12049_/X
+ sky130_fd_sc_hd__o211a_1
X_16926_ _17870_/CLK _16926_/D vssd1 vssd1 vccd1 vccd1 _16926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16857_ _18060_/CLK _16857_/D vssd1 vssd1 vccd1 vccd1 _16857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15808_ _17725_/CLK _15808_/D vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16788_ _18055_/CLK _16788_/D vssd1 vssd1 vccd1 vccd1 _16788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15739_ _17742_/CLK _15739_/D vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09260_ _12756_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _16241_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18458_ _18458_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08211_ _15545_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17409_ _17439_/CLK _17409_/D vssd1 vssd1 vccd1 vccd1 _17409_/Q sky130_fd_sc_hd__dfxtp_1
X_09191_ hold2376/X _09216_/B _09190_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _09191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18389_ _18389_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08142_ hold173/X _15710_/Q hold196/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__mux2_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08073_ hold1049/X _08082_/B _08072_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _08073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4003 _16540_/Q vssd1 vssd1 vccd1 vccd1 hold4003/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4014 _16435_/Q vssd1 vssd1 vccd1 vccd1 hold4014/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4025 _12004_/X vssd1 vssd1 vccd1 vccd1 _17158_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4036 _10723_/X vssd1 vssd1 vccd1 vccd1 _16731_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3302 _12926_/X vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4047 _16473_/Q vssd1 vssd1 vccd1 vccd1 hold4047/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4058 _10417_/X vssd1 vssd1 vccd1 vccd1 _16629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3313 _17591_/Q vssd1 vssd1 vccd1 vccd1 hold3313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3324 _17718_/Q vssd1 vssd1 vccd1 vccd1 hold3324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4069 _17654_/Q vssd1 vssd1 vccd1 vccd1 hold4069/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3335 _10201_/X vssd1 vssd1 vccd1 vccd1 _16557_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3346 _17380_/Q vssd1 vssd1 vccd1 vccd1 hold3346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2601 _17955_/Q vssd1 vssd1 vccd1 vccd1 hold2601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2612 _18168_/Q vssd1 vssd1 vccd1 vccd1 hold2612/X sky130_fd_sc_hd__dlygate4sd3_1
X_08975_ hold5/X hold329/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__mux2_1
Xhold3357 _17632_/Q vssd1 vssd1 vccd1 vccd1 hold3357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 _07905_/X vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3368 _17237_/Q vssd1 vssd1 vccd1 vccd1 hold3368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__buf_4
Xhold3379 _09646_/X vssd1 vssd1 vccd1 vccd1 _16372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _14973_/X vssd1 vssd1 vccd1 vccd1 _18272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 _09292_/X vssd1 vssd1 vccd1 vccd1 _16256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1900 _14911_/X vssd1 vssd1 vccd1 vccd1 _18243_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _15549_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__or2_1
Xhold2656 _16278_/Q vssd1 vssd1 vccd1 vccd1 hold2656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 _18070_/Q vssd1 vssd1 vccd1 vccd1 hold1911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 la_data_in[27] vssd1 vssd1 vccd1 vccd1 hold581/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2667 _14121_/X vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__buf_4
Xhold1933 _14899_/X vssd1 vssd1 vccd1 vccd1 _18237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 _16251_/Q vssd1 vssd1 vccd1 vccd1 hold2678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _15636_/Q vssd1 vssd1 vccd1 vccd1 hold2689/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1944 _07977_/X vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 _07961_/X vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1966 _15578_/Q vssd1 vssd1 vccd1 vccd1 hold1966/X sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _14529_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07857_/X sky130_fd_sc_hd__or2_1
Xhold1977 _17907_/Q vssd1 vssd1 vccd1 vccd1 hold1977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1988 _08271_/X vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1999 _14089_/X vssd1 vssd1 vccd1 vccd1 _17849_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07788_ _07788_/A vssd1 vssd1 vccd1 vccd1 _07788_/Y sky130_fd_sc_hd__inv_2
X_09527_ hold2497/X _16333_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09463_/C _09463_/D _09481_/B vssd1 vssd1 vccd1 vccd1 _09458_/Y sky130_fd_sc_hd__a21boi_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ hold949/X _08445_/B vssd1 vssd1 vccd1 vccd1 _08409_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _07805_/A _09362_/A _09362_/D vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__a21o_1
X_11420_ hold2505/X hold3392/X _11741_/C vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11351_ hold2597/X _16941_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10302_ _10542_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ _14517_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11282_ hold2877/X hold5324/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__mux2_1
Xhold5260 _16732_/Q vssd1 vssd1 vccd1 vccd1 hold5260/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_13021_ _13048_/A hold900/X hold616/X vssd1 vssd1 vccd1 vccd1 hold901/A sky130_fd_sc_hd__a21o_1
Xhold5271 _10027_/Y vssd1 vssd1 vccd1 vccd1 _16499_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _10548_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__or2_1
Xhold5282 _11751_/Y vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5293 _10030_/Y vssd1 vssd1 vccd1 vccd1 _16500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4570 _11845_/X vssd1 vssd1 vccd1 vccd1 _17105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4581 _16700_/Q vssd1 vssd1 vccd1 vccd1 hold4581/X sky130_fd_sc_hd__dlygate4sd3_1
X_10164_ _10548_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__or2_1
Xhold4592 _10708_/X vssd1 vssd1 vccd1 vccd1 _16726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3880 _17101_/Q vssd1 vssd1 vccd1 vccd1 hold3880/X sky130_fd_sc_hd__dlygate4sd3_1
X_14972_ _14972_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or2_1
Xhold3891 _11485_/X vssd1 vssd1 vccd1 vccd1 _16985_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17760_ _17855_/CLK _17760_/D vssd1 vssd1 vccd1 vccd1 _17760_/Q sky130_fd_sc_hd__dfxtp_1
X_10095_ _11082_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__or2_1
X_13923_ _13923_/A hold736/X vssd1 vssd1 vccd1 vccd1 hold737/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16711_ _18042_/CLK _16711_/D vssd1 vssd1 vccd1 vccd1 _16711_/Q sky130_fd_sc_hd__dfxtp_1
X_17691_ _17691_/CLK _17691_/D vssd1 vssd1 vccd1 vccd1 _17691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16642_ _18224_/CLK _16642_/D vssd1 vssd1 vccd1 vccd1 _16642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ hold4169/X _13788_/A _13853_/X vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ hold2520/X _17446_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__mux2_1
X_16573_ _18131_/CLK _16573_/D vssd1 vssd1 vccd1 vccd1 _16573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _13788_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13785_/X sky130_fd_sc_hd__or2_1
X_10997_ hold1569/X _16823_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__mux2_1
X_18312_ _18373_/CLK hold267/X vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_15524_ hold1014/X _15560_/A2 _15523_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _15524_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ hold917/X hold3038/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18243_ _18243_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15455_ _15455_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__or2_1
X_12667_ hold2062/X hold2864/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14406_ hold2947/X hold209/X _14405_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _14406_/X
+ sky130_fd_sc_hd__o211a_1
X_18174_ _18206_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
X_11618_ hold2060/X hold4881/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__mux2_1
X_15386_ _17342_/Q _09362_/C _09362_/D hold674/X vssd1 vssd1 vccd1 vccd1 _15386_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ hold1311/X hold3008/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _17260_/CLK _17125_/D vssd1 vssd1 vccd1 vccd1 _17125_/Q sky130_fd_sc_hd__dfxtp_1
X_14337_ hold2917/X _14326_/B _14336_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14337_/X
+ sky130_fd_sc_hd__o211a_1
X_11549_ hold2236/X _17007_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__mux2_1
Xhold507 hold507/A vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 hold518/A vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold529 hold529/A vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ _17893_/CLK _17056_/D vssd1 vssd1 vccd1 vccd1 _17056_/Q sky130_fd_sc_hd__dfxtp_1
X_14268_ _15217_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16007_ _18414_/CLK _16007_/D vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
X_13219_ _13218_/X hold5898/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ hold2230/X _14198_/B _14198_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _14199_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _07943_/X vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _15314_/A _08760_/B vssd1 vssd1 vccd1 vccd1 _16000_/D sky130_fd_sc_hd__and2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _15739_/Q vssd1 vssd1 vccd1 vccd1 hold1218/X sky130_fd_sc_hd__dlygate4sd3_1
X_17958_ _18208_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_81_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1229 _17782_/Q vssd1 vssd1 vccd1 vccd1 hold1229/X sky130_fd_sc_hd__dlygate4sd3_1
X_16909_ _17856_/CLK _16909_/D vssd1 vssd1 vccd1 vccd1 _16909_/Q sky130_fd_sc_hd__dfxtp_1
X_08691_ hold59/X hold701/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08692_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17889_ _17889_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ hold2951/X _09325_/B _09311_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09312_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ _15519_/A hold2238/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _15557_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _13939_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _15701_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ _15515_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08056_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3110 _12875_/X vssd1 vssd1 vccd1 vccd1 _12876_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3121 _17476_/Q vssd1 vssd1 vccd1 vccd1 hold3121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3132 _16532_/Q vssd1 vssd1 vccd1 vccd1 hold3132/X sky130_fd_sc_hd__buf_1
Xhold3143 _12310_/Y vssd1 vssd1 vccd1 vccd1 _17260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3154 _12351_/Y vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2420 _14773_/X vssd1 vssd1 vccd1 vccd1 _18177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3165 _17095_/Q vssd1 vssd1 vccd1 vccd1 hold3165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2431 _15828_/Q vssd1 vssd1 vccd1 vccd1 hold2431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3176 _12334_/Y vssd1 vssd1 vccd1 vccd1 _17268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08958_ _15473_/A hold305/X vssd1 vssd1 vccd1 vccd1 _16096_/D sky130_fd_sc_hd__and2_1
Xhold3187 _13888_/Y vssd1 vssd1 vccd1 vccd1 _17749_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2442 _08042_/X vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2453 _18121_/Q vssd1 vssd1 vccd1 vccd1 hold2453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3198 _13849_/Y vssd1 vssd1 vccd1 vccd1 _17736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2464 _15799_/Q vssd1 vssd1 vccd1 vccd1 hold2464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 _13038_/X vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2475 _15719_/Q vssd1 vssd1 vccd1 vccd1 hold2475/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1741 _08077_/X vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07909_ hold1134/X _07918_/B _07908_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07909_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2486 _14255_/X vssd1 vssd1 vccd1 vccd1 _17928_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _16162_/Q vssd1 vssd1 vccd1 vccd1 hold1752/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2497 _18246_/Q vssd1 vssd1 vccd1 vccd1 hold2497/X sky130_fd_sc_hd__dlygate4sd3_1
X_08889_ _13002_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _16062_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1763 _18361_/Q vssd1 vssd1 vccd1 vccd1 hold1763/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 _07825_/X vssd1 vssd1 vccd1 vccd1 _17751_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _11031_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__or2_1
Xhold1785 _14569_/X vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1796 _14563_/X vssd1 vssd1 vccd1 vccd1 _18076_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10851_ _11616_/A _10851_/B vssd1 vssd1 vccd1 vccd1 _10851_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ hold4641/X _13856_/B _13569_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13570_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _11106_/A _10782_/B vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__or2_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ hold3046/X _12520_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__mux2_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15240_ hold89/X _15486_/A2 _15446_/B1 _16053_/Q vssd1 vssd1 vccd1 vccd1 _15240_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _17319_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _12234_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15171_ hold573/X _15179_/B vssd1 vssd1 vccd1 vccd1 _15171_/X sky130_fd_sc_hd__or2_1
X_12383_ hold68/X hold473/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12384_/B sky130_fd_sc_hd__mux2_1
X_14122_ _14246_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14122_/X sky130_fd_sc_hd__or2_1
X_11334_ _12204_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ hold2163/X _14036_/B _14052_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14053_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _12093_/A _11265_/B vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or2_1
Xhold5090 _17084_/Q vssd1 vssd1 vccd1 vccd1 hold5090/X sky130_fd_sc_hd__dlygate4sd3_1
X_13004_ _14897_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _13017_/B sky130_fd_sc_hd__or2_2
X_10216_ hold3965/X _10643_/B _10215_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ hold5263/X _11115_/A _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17812_ _18427_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_1
X_10147_ hold3976/X _10643_/B _10146_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14955_ hold861/X _14946_/B _14954_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 hold862/A
+ sky130_fd_sc_hd__o211a_1
X_17743_ _17743_/CLK _17743_/D vssd1 vssd1 vccd1 vccd1 _17743_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ hold5116/X _11192_/B _10077_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10078_/X
+ sky130_fd_sc_hd__o211a_1
X_13906_ _14246_/A hold2850/X hold244/X vssd1 vssd1 vccd1 vccd1 _13907_/B sky130_fd_sc_hd__mux2_1
X_14886_ _15225_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14886_/X sky130_fd_sc_hd__or2_1
X_17674_ _17738_/CLK _17674_/D vssd1 vssd1 vccd1 vccd1 _17674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16625_ _18131_/CLK _16625_/D vssd1 vssd1 vccd1 vccd1 _16625_/Q sky130_fd_sc_hd__dfxtp_1
X_13837_ _13873_/A _13837_/B vssd1 vssd1 vccd1 vccd1 _13837_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _18210_/CLK _16556_/D vssd1 vssd1 vccd1 vccd1 _16556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13768_ hold3277/X _13862_/B _13767_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13768_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12719_ hold3489/X _12718_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__mux2_1
X_15507_ _15508_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _15507_/Y sky130_fd_sc_hd__nor2_1
X_16487_ _18415_/CLK _16487_/D vssd1 vssd1 vccd1 vccd1 _16487_/Q sky130_fd_sc_hd__dfxtp_1
X_13699_ hold3324/X _13829_/B _13698_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13699_/X
+ sky130_fd_sc_hd__o211a_1
X_15438_ hold268/X _09367_/A _15486_/B1 _17347_/Q vssd1 vssd1 vccd1 vccd1 _15438_/X
+ sky130_fd_sc_hd__a22o_1
X_18226_ _18226_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18157_ _18221_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
X_15369_ hold590/X _15485_/A2 _15447_/B1 hold470/X _15368_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17108_ _17268_/CLK _17108_/D vssd1 vssd1 vccd1 vccd1 _17108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold315 input33/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18088_ _18126_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 hold337/A vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _09948_/A _09930_/B vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__or2_1
X_17039_ _17887_/CLK _17039_/D vssd1 vssd1 vccd1 vccd1 _17039_/Q sky130_fd_sc_hd__dfxtp_1
Xhold359 hold29/X vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 _15208_/C1 vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__buf_4
XFILLER_0_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09861_ _09933_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout817 _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14879_/C1 sky130_fd_sc_hd__buf_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 fanout841/X vssd1 vssd1 vccd1 vccd1 _14807_/C1 sky130_fd_sc_hd__buf_4
Xfanout839 _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14877_/C1 sky130_fd_sc_hd__buf_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ hold32/X hold673/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _18390_/Q vssd1 vssd1 vccd1 vccd1 hold1004/X sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ _09987_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__or2_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _15524_/X vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _08118_/X vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ hold26/X hold597/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__mux2_1
Xhold1037 la_data_in[11] vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _14129_/X vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _14794_/X vssd1 vssd1 vccd1 vccd1 hold1059/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _15454_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _15958_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_287_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_216_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18069_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ hold800/X _09230_/B vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ hold1185/X _09177_/A2 _09156_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _15513_/A hold2994/X hold196/X vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ _14988_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _14726_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08039_/X sky130_fd_sc_hd__or2_1
Xhold860 hold860/A vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 hold871/A vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 hold882/A vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 hold893/A vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ hold4659/X _11732_/B _11049_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11050_/X
+ sky130_fd_sc_hd__o211a_1
X_10001_ _16491_/Q _10001_/B _10001_/C vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__and3_1
XFILLER_0_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 _16165_/Q vssd1 vssd1 vccd1 vccd1 hold2250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2261 _07903_/X vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2272 _18280_/Q vssd1 vssd1 vccd1 vccd1 hold2272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2283 _18221_/Q vssd1 vssd1 vccd1 vccd1 hold2283/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _14731_/X vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _14871_/X vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1571 _18251_/Q vssd1 vssd1 vccd1 vccd1 hold1571/X sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ _14740_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__or2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _12153_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__or2_1
Xhold1582 _18232_/Q vssd1 vssd1 vccd1 vccd1 hold1582/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1593 _18217_/Q vssd1 vssd1 vccd1 vccd1 hold1593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ hold5346/X _11216_/B _10902_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _10903_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ hold1440/X _14666_/B _14670_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14671_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _13392_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _18355_/CLK _16410_/D vssd1 vssd1 vccd1 vccd1 _16410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13622_ hold1822/X _17661_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__mux2_1
X_17390_ _18451_/CLK _17390_/D vssd1 vssd1 vccd1 vccd1 _17390_/Q sky130_fd_sc_hd__dfxtp_1
X_10834_ hold5518/X _11216_/B _10833_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10834_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _18382_/CLK _16341_/D vssd1 vssd1 vccd1 vccd1 _16341_/Q sky130_fd_sc_hd__dfxtp_1
X_13553_ hold1024/X hold4826/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ hold3240/X _11156_/B _10764_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10765_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12504_ _17345_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__or2_1
X_16272_ _17375_/CLK _16272_/D vssd1 vssd1 vccd1 vccd1 _16272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13484_ hold1513/X _17615_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__mux2_1
X_10696_ hold5488/X _11210_/B _10695_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _10696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15223_ hold730/X _15233_/B vssd1 vssd1 vccd1 vccd1 _15223_/X sky130_fd_sc_hd__or2_1
X_18011_ _18431_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
X_12435_ hold44/X hold222/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12436_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ hold1663/X _15161_/B _15153_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o211a_1
X_12366_ hold3162/X _12279_/A _12365_/X vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ hold1434/X _14105_/A2 _14104_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14105_/X
+ sky130_fd_sc_hd__o211a_1
X_11317_ hold5064/X _12341_/B _11316_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11317_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15085_ _15193_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__or2_1
X_12297_ hold3775/X _13716_/A _12296_/X vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__a21oi_1
X_14036_ _15543_/A _14036_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ hold4617/X _11726_/B _11247_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11248_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _11194_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11179_/Y sky130_fd_sc_hd__nor2_1
X_15987_ _18414_/CLK _15987_/D vssd1 vssd1 vccd1 vccd1 hold401/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17726_ _17726_/CLK _17726_/D vssd1 vssd1 vccd1 vccd1 _17726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14938_ _15207_/A _14962_/B vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _17721_/CLK _17657_/D vssd1 vssd1 vccd1 vccd1 _17657_/Q sky130_fd_sc_hd__dfxtp_1
X_14869_ hold2891/X _14880_/B _14868_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16608_ _18225_/CLK _16608_/D vssd1 vssd1 vccd1 vccd1 _16608_/Q sky130_fd_sc_hd__dfxtp_1
X_08390_ _14786_/A hold2108/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__mux2_1
X_17588_ _17715_/CLK _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _18225_/CLK _16539_/D vssd1 vssd1 vccd1 vccd1 _16539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _16122_/D sky130_fd_sc_hd__and2_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18209_ _18268_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5804 hold5929/X vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5815 _18411_/Q vssd1 vssd1 vccd1 vccd1 hold5815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 input18/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__buf_1
Xhold5826 _18402_/Q vssd1 vssd1 vccd1 vccd1 hold5826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5837 _17522_/Q vssd1 vssd1 vccd1 vccd1 hold5837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5848 hold5940/X vssd1 vssd1 vccd1 vccd1 hold5848/X sky130_fd_sc_hd__clkbuf_2
Xhold134 hold1/X vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5859 hold5859/A vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_12
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 input11/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ hold5429/X _10025_/B _09912_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _09484_/B vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout614 _09358_/Y vssd1 vssd1 vccd1 vccd1 _15487_/B1 sky130_fd_sc_hd__buf_6
Xfanout625 _09347_/Y vssd1 vssd1 vccd1 vccd1 _15484_/A2 sky130_fd_sc_hd__buf_6
Xfanout636 fanout660/X vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__clkbuf_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout647 _12885_/A vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__buf_4
X_09844_ hold5745/X _10016_/B _09843_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09844_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout658 _14360_/A vssd1 vssd1 vccd1 vccd1 _15504_/A sky130_fd_sc_hd__buf_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 _08137_/A vssd1 vssd1 vccd1 vccd1 _13723_/C1 sky130_fd_sc_hd__buf_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ hold3491/X _10073_/B _09774_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09775_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _15050_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _15984_/D sky130_fd_sc_hd__and2_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ hold380/X hold699/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__mux2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08588_ hold359/X hold553/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ hold1582/X _16674_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09209_ hold2365/X _09218_/B _09208_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _09209_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10481_ hold1337/X _16651_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12220_ _12314_/A _12314_/B _12219_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ hold4723/X _12377_/B _12150_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ hold1727/X hold5536/X _11213_/C vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12082_ hold3372/X _12374_/B _12081_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _17184_/D
+ sky130_fd_sc_hd__o211a_1
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
X_15910_ _17307_/CLK _15910_/D vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__dfxtp_1
X_11033_ hold2068/X hold5661/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__mux2_1
X_16890_ _18061_/CLK _16890_/D vssd1 vssd1 vccd1 vccd1 _16890_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _17732_/CLK _15841_/D vssd1 vssd1 vccd1 vccd1 _15841_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _17938_/Q vssd1 vssd1 vccd1 vccd1 hold2080/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18392_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2091 _15744_/Q vssd1 vssd1 vccd1 vccd1 hold2091/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _17691_/CLK _15772_/D vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfxtp_1
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _17504_/D sky130_fd_sc_hd__and2_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 _14993_/X vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17511_/CLK _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
X_14723_ hold1952/X _14718_/B _14722_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14723_/X
+ sky130_fd_sc_hd__o211a_1
X_11935_ hold5026/X _12356_/B _11934_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14654_ _15209_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14654_/X sky130_fd_sc_hd__or2_1
X_17442_ _17448_/CLK _17442_/D vssd1 vssd1 vccd1 vccd1 _17442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ hold3362/X _13844_/B _11865_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11866_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13800_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ hold1936/X hold4035/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17373_ _17375_/CLK _17373_/D vssd1 vssd1 vccd1 vccd1 _17373_/Q sky130_fd_sc_hd__dfxtp_1
X_14585_ hold2999/X _14612_/B _14584_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ _12343_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ _13737_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16324_ _18397_/CLK _16324_/D vssd1 vssd1 vccd1 vccd1 _16324_/Q sky130_fd_sc_hd__dfxtp_1
X_10748_ _17943_/Q hold3202/X _11735_/C vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _17487_/CLK _16255_/D vssd1 vssd1 vccd1 vccd1 _16255_/Q sky130_fd_sc_hd__dfxtp_1
X_13467_ _13788_/A _13467_/B vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__or2_1
X_10679_ hold2699/X hold3665/X _11735_/C vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15206_ hold2748/X _15221_/B _15205_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15206_/X
+ sky130_fd_sc_hd__o211a_1
X_12418_ _12420_/A hold547/X vssd1 vssd1 vccd1 vccd1 _17302_/D sky130_fd_sc_hd__and2_1
X_16186_ _17482_/CLK _16186_/D vssd1 vssd1 vccd1 vccd1 _16186_/Q sky130_fd_sc_hd__dfxtp_1
X_13398_ _13791_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _15191_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _13873_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3709 _11193_/Y vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__dlygate4sd3_1
X_15068_ _15068_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__and2_1
X_14019_ hold2620/X _14040_/B _14018_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14019_/X
+ sky130_fd_sc_hd__o211a_1
X_07890_ _14740_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07890_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ hold1671/X _13222_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__mux2_1
X_08511_ _15515_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__or2_1
X_17709_ _17741_/CLK _17709_/D vssd1 vssd1 vccd1 vccd1 _17709_/Q sky130_fd_sc_hd__dfxtp_1
X_09491_ _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13056_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_176_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ hold2401/X _08433_/B _08441_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08442_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_25__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_25__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ _08373_/A hold123/X vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__and2_1
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5601 _09805_/X vssd1 vssd1 vccd1 vccd1 _16425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5612 _16423_/Q vssd1 vssd1 vccd1 vccd1 hold5612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5623 _16869_/Q vssd1 vssd1 vccd1 vccd1 hold5623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5634 _11272_/X vssd1 vssd1 vccd1 vccd1 _16914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4900 _12031_/X vssd1 vssd1 vccd1 vccd1 _17167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5645 _16886_/Q vssd1 vssd1 vccd1 vccd1 hold5645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4911 _16968_/Q vssd1 vssd1 vccd1 vccd1 hold4911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5656 _09502_/X vssd1 vssd1 vccd1 vccd1 _16324_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5667 _09640_/X vssd1 vssd1 vccd1 vccd1 _16370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4922 _10852_/X vssd1 vssd1 vccd1 vccd1 _16774_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4933 _17272_/Q vssd1 vssd1 vccd1 vccd1 hold4933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5678 _11311_/X vssd1 vssd1 vccd1 vccd1 _16927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4944 _13759_/X vssd1 vssd1 vccd1 vccd1 _17706_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5689 _17078_/Q vssd1 vssd1 vccd1 vccd1 hold5689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4955 _17615_/Q vssd1 vssd1 vccd1 vccd1 hold4955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4966 _12025_/X vssd1 vssd1 vccd1 vccd1 _17165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout400 _14447_/Y vssd1 vssd1 vccd1 vccd1 _14481_/B sky130_fd_sc_hd__clkbuf_8
Xhold4977 _16648_/Q vssd1 vssd1 vccd1 vccd1 hold4977/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout411 _14232_/Y vssd1 vssd1 vccd1 vccd1 _14266_/B sky130_fd_sc_hd__buf_6
Xfanout422 _14036_/B vssd1 vssd1 vccd1 vccd1 _14040_/B sky130_fd_sc_hd__clkbuf_8
Xhold4988 _11140_/X vssd1 vssd1 vccd1 vccd1 _16870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4999 _16471_/Q vssd1 vssd1 vccd1 vccd1 hold4999/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout433 _13052_/X vssd1 vssd1 vccd1 vccd1 _13183_/A1 sky130_fd_sc_hd__buf_6
Xfanout444 _12353_/C vssd1 vssd1 vccd1 vccd1 _13793_/S sky130_fd_sc_hd__clkbuf_8
Xfanout455 _11171_/C vssd1 vssd1 vccd1 vccd1 _11735_/C sky130_fd_sc_hd__clkbuf_8
Xfanout466 _13886_/C vssd1 vssd1 vccd1 vccd1 _13880_/C sky130_fd_sc_hd__clkbuf_8
X_09827_ hold1332/X hold5379/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__mux2_1
Xfanout477 _11672_/S vssd1 vssd1 vccd1 vccd1 _12152_/S sky130_fd_sc_hd__clkbuf_8
Xfanout488 _10874_/S vssd1 vssd1 vccd1 vccd1 _11201_/C sky130_fd_sc_hd__clkbuf_8
Xfanout499 _10562_/S vssd1 vssd1 vccd1 vccd1 _11192_/C sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_231_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17279_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ hold1690/X _16410_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__mux2_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08709_ hold140/X hold530/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__mux2_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ hold1656/X hold5134/X _10481_/S vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _17064_/Q _12299_/B _12299_/C vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__and3_1
XFILLER_0_178_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ hold1043/X _17041_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__mux2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10602_ hold3179/X _10098_/A _10601_/X vssd1 vssd1 vccd1 vccd1 _10602_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14370_ _14376_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _17984_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11582_ hold1309/X _17018_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ hold3217/X _13814_/B _13320_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__o211a_1
X_10533_ _10551_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16040_ _18423_/CLK _16040_/D vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13252_ hold5260/X _13251_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__mux2_2
X_10464_ _10560_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ hold2316/X hold4655/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _13183_/A1 _13181_/X _13182_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13183_/X
+ sky130_fd_sc_hd__o211a_1
X_10395_ _10527_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ hold2133/X _17202_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__mux2_1
X_17991_ _18055_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_319_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12065_ hold2963/X hold4712/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__mux2_1
X_16942_ _18051_/CLK _16942_/D vssd1 vssd1 vccd1 vccd1 _16942_/Q sky130_fd_sc_hd__dfxtp_1
X_11016_ _11031_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__or2_1
X_16873_ _18013_/CLK _16873_/D vssd1 vssd1 vccd1 vccd1 _16873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _17738_/CLK _15824_/D vssd1 vssd1 vccd1 vccd1 _15824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _17740_/CLK _15755_/D vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfxtp_1
X_12967_ hold2582/X hold3057/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__mux2_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _15099_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__or2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ hold2185/X hold3320/X _13811_/C vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__mux2_1
X_15686_ _17274_/CLK _15686_/D vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfxtp_1
X_12898_ hold1975/X hold3004/X _12910_/S vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17425_ _17629_/CLK _17425_/D vssd1 vssd1 vccd1 vccd1 _17425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14637_ hold1723/X _14666_/B _14636_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14637_/X
+ sky130_fd_sc_hd__o211a_1
X_11849_ hold2468/X hold5239/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11850_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17356_ _17487_/CLK _17356_/D vssd1 vssd1 vccd1 vccd1 _17356_/Q sky130_fd_sc_hd__dfxtp_1
X_14568_ _15492_/A _14573_/B hold1783/X vssd1 vssd1 vccd1 vccd1 _14568_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18073_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16307_ _17511_/CLK _16307_/D vssd1 vssd1 vccd1 vccd1 _16307_/Q sky130_fd_sc_hd__dfxtp_1
X_13519_ hold3251/X _13808_/B _13518_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13519_/X
+ sky130_fd_sc_hd__o211a_1
X_17287_ _17287_/CLK _17287_/D vssd1 vssd1 vccd1 vccd1 hold594/A sky130_fd_sc_hd__dfxtp_1
X_14499_ hold784/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16238_ _17419_/CLK _16238_/D vssd1 vssd1 vccd1 vccd1 _16238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4207 _17727_/Q vssd1 vssd1 vccd1 vccd1 hold4207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4218 _17162_/Q vssd1 vssd1 vccd1 vccd1 hold4218/X sky130_fd_sc_hd__dlygate4sd3_1
X_16169_ _17503_/CLK _16169_/D vssd1 vssd1 vccd1 vccd1 _16169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4229 _10984_/X vssd1 vssd1 vccd1 vccd1 _16818_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3506 _17449_/Q vssd1 vssd1 vccd1 vccd1 hold3506/X sky130_fd_sc_hd__dlygate4sd3_1
X_08991_ hold359/X hold361/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__mux2_1
Xhold3517 _17446_/Q vssd1 vssd1 vccd1 vccd1 hold3517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3528 _17441_/Q vssd1 vssd1 vccd1 vccd1 hold3528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3539 _17717_/Q vssd1 vssd1 vccd1 vccd1 hold3539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2805 _15671_/Q vssd1 vssd1 vccd1 vccd1 hold2805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2816 _18333_/Q vssd1 vssd1 vccd1 vccd1 hold2816/X sky130_fd_sc_hd__dlygate4sd3_1
X_07942_ hold756/X _07988_/B vssd1 vssd1 vccd1 vccd1 _07942_/X sky130_fd_sc_hd__or2_1
Xhold2827 _09081_/X vssd1 vssd1 vccd1 vccd1 _16155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_9__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_9__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
Xhold2838 _18276_/Q vssd1 vssd1 vccd1 vccd1 hold2838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2849 _14526_/X vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07873_ _14330_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ _09903_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09612_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09543_ _09987_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09474_ hold681/X _09477_/C _09481_/B vssd1 vssd1 vccd1 vccd1 _09474_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08425_ _15539_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _15525_/A hold2561/X hold122/X vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ hold756/X _08335_/B vssd1 vssd1 vccd1 vccd1 _08287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5420 _09823_/X vssd1 vssd1 vccd1 vccd1 _16431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5431 _16885_/Q vssd1 vssd1 vccd1 vccd1 hold5431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5442 _11080_/X vssd1 vssd1 vccd1 vccd1 _16850_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5453 _10735_/X vssd1 vssd1 vccd1 vccd1 _16735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5464 _16894_/Q vssd1 vssd1 vccd1 vccd1 hold5464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4730 _12094_/X vssd1 vssd1 vccd1 vccd1 _17188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5475 _11119_/X vssd1 vssd1 vccd1 vccd1 _16863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4741 hold5829/X vssd1 vssd1 vccd1 vccd1 hold5830/A sky130_fd_sc_hd__buf_4
Xhold5486 _16990_/Q vssd1 vssd1 vccd1 vccd1 hold5486/X sky130_fd_sc_hd__dlygate4sd3_1
X_10180_ hold4698/X _10568_/B _10179_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10180_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4752 _10840_/X vssd1 vssd1 vccd1 vccd1 _16770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5497 _09802_/X vssd1 vssd1 vccd1 vccd1 _16424_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4763 _17155_/Q vssd1 vssd1 vccd1 vccd1 hold4763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4774 _12268_/X vssd1 vssd1 vccd1 vccd1 _17246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4785 _17231_/Q vssd1 vssd1 vccd1 vccd1 hold4785/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout230 _10610_/B vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__buf_4
Xhold4796 _11863_/X vssd1 vssd1 vccd1 vccd1 _17111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout241 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _09952_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _12210_/A vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__buf_4
Xfanout263 _11616_/A vssd1 vssd1 vccd1 vccd1 _12018_/A sky130_fd_sc_hd__buf_4
Xfanout274 _13770_/A vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__clkbuf_4
Xfanout285 fanout298/X vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__clkbuf_4
Xfanout296 _11031_/A vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__buf_4
X_13870_ _13873_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nor2_1
X_12821_ hold3469/X _12820_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12752_ hold3025/X _12751_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__mux2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ hold1480/X _15547_/B _15539_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ _12153_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__or2_1
X_15471_ _15471_/A _15471_/B _15471_/C _15471_/D vssd1 vssd1 vccd1 vccd1 _15471_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ hold3089/X _12682_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17274_/CLK _17210_/D vssd1 vssd1 vccd1 vccd1 _17210_/Q sky130_fd_sc_hd__dfxtp_1
X_14422_ hold1778/X _14433_/B _14421_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _14422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11634_ _11637_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__or2_1
X_18190_ _18190_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17141_ _17208_/CLK _17141_/D vssd1 vssd1 vccd1 vccd1 _17141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14980_/A hold2853/X hold275/X vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11565_ _11667_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__or2_1
X_13304_ _13297_/X _13303_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__o21a_1
X_10516_ hold4263/X _10610_/B _10515_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10516_/X
+ sky130_fd_sc_hd__o211a_1
X_17072_ _18427_/CLK _17072_/D vssd1 vssd1 vccd1 vccd1 _17072_/Q sky130_fd_sc_hd__dfxtp_1
X_14284_ hold784/X _14284_/B vssd1 vssd1 vccd1 vccd1 hold785/A sky130_fd_sc_hd__or2_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11496_ _11688_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11496_/X sky130_fd_sc_hd__or2_1
X_16023_ _17530_/CLK _16023_/D vssd1 vssd1 vccd1 vccd1 hold660/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13235_ _13234_/X _16922_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__mux2_1
X_10447_ hold3271/X _10631_/B _10446_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ _13166_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__or2_1
X_10378_ hold4977/X _10628_/B _10377_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_153_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18229_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12117_ _13797_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13097_ _13097_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__and2_1
X_17974_ _18069_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
X_12048_ _12282_/A _12048_/B vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__or2_1
X_16925_ _17901_/CLK _16925_/D vssd1 vssd1 vccd1 vccd1 _16925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16856_ _18059_/CLK _16856_/D vssd1 vssd1 vccd1 vccd1 _16856_/Q sky130_fd_sc_hd__dfxtp_1
X_15807_ _17686_/CLK _15807_/D vssd1 vssd1 vccd1 vccd1 _15807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16787_ _18054_/CLK _16787_/D vssd1 vssd1 vccd1 vccd1 _16787_/Q sky130_fd_sc_hd__dfxtp_1
X_13999_ hold2026/X _13986_/B _13998_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 _13999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _17741_/CLK _15738_/D vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18457_ _18458_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ _17878_/CLK _15669_/D vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ hold2032/X _08209_/B _08209_/Y _08141_/A vssd1 vssd1 vccd1 vccd1 _08210_/X
+ sky130_fd_sc_hd__o211a_1
X_17408_ _18458_/CLK _17408_/D vssd1 vssd1 vccd1 vccd1 _17408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _15519_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__or2_1
X_18388_ _18388_/CLK hold988/X vssd1 vssd1 vccd1 vccd1 hold987/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08141_ _08141_/A hold517/X vssd1 vssd1 vccd1 vccd1 _15709_/D sky130_fd_sc_hd__and2_1
X_17339_ _17343_/CLK hold57/X vssd1 vssd1 vccd1 vccd1 _17339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _14866_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4004 _10629_/Y vssd1 vssd1 vccd1 vccd1 _10630_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4015 _09739_/X vssd1 vssd1 vccd1 vccd1 _16403_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4026 _16871_/Q vssd1 vssd1 vccd1 vccd1 hold4026/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4037 hold5840/X vssd1 vssd1 vccd1 vccd1 hold5841/A sky130_fd_sc_hd__buf_4
Xhold4048 _09853_/X vssd1 vssd1 vccd1 vccd1 _16441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3303 _17462_/Q vssd1 vssd1 vccd1 vccd1 hold3303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4059 _16467_/Q vssd1 vssd1 vccd1 vccd1 hold4059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3314 _13318_/X vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3325 _13699_/X vssd1 vssd1 vccd1 vccd1 _17686_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3336 _17600_/Q vssd1 vssd1 vccd1 vccd1 hold3336/X sky130_fd_sc_hd__dlygate4sd3_1
X_08974_ _12428_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _16104_/D sky130_fd_sc_hd__and2_1
Xhold3347 _17184_/Q vssd1 vssd1 vccd1 vccd1 hold3347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2602 _14311_/X vssd1 vssd1 vccd1 vccd1 _17955_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3358 _16509_/Q vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _14755_/X vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2624 _16208_/Q vssd1 vssd1 vccd1 vccd1 hold2624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3369 _12145_/X vssd1 vssd1 vccd1 vccd1 _17205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold73/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _16159_/Q vssd1 vssd1 vccd1 vccd1 hold2635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ hold1792/X _07924_/B _07924_/Y _08161_/A vssd1 vssd1 vccd1 vccd1 _07925_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1901 _15655_/Q vssd1 vssd1 vccd1 vccd1 hold1901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_2
Xhold2646 _15667_/Q vssd1 vssd1 vccd1 vccd1 hold2646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 _09336_/X vssd1 vssd1 vccd1 vccd1 _16278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 _14548_/X vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _16194_/Q vssd1 vssd1 vccd1 vccd1 hold1923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _18176_/Q vssd1 vssd1 vccd1 vccd1 hold2668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _15796_/Q vssd1 vssd1 vccd1 vccd1 hold1934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 _15804_/Q vssd1 vssd1 vccd1 vccd1 hold2679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1945 _16218_/Q vssd1 vssd1 vccd1 vccd1 hold1945/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ hold2687/X _07869_/B _07855_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07856_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1956 _17911_/Q vssd1 vssd1 vccd1 vccd1 hold1956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1967 _07866_/X vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 _14209_/X vssd1 vssd1 vccd1 vccd1 _17907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _17995_/Q vssd1 vssd1 vccd1 vccd1 hold1989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07787_ _12343_/A vssd1 vssd1 vccd1 vccd1 _07787_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_151_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ hold5338/X _10013_/B _09525_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09463_/D _09481_/B _09457_/C vssd1 vssd1 vccd1 vccd1 _16312_/D sky130_fd_sc_hd__and3b_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ hold2546/X _08440_/A2 _08407_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ hold5851/A _09342_/B _09342_/Y _09387_/X _12442_/A vssd1 vssd1 vccd1 vccd1
+ _09388_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08339_ _08504_/A hold300/A vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ hold3537/X _11617_/A2 _11349_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ hold2070/X _16591_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__mux2_1
X_11281_ hold5737/X _11765_/B _11280_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ _09489_/B hold927/A vssd1 vssd1 vccd1 vccd1 hold900/A sky130_fd_sc_hd__nand2b_1
Xhold5250 _11218_/Y vssd1 vssd1 vccd1 vccd1 _16896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5261 _11205_/Y vssd1 vssd1 vccd1 vccd1 _11206_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10232_ hold2359/X _16568_/Q _10643_/C vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5272 _16926_/Q vssd1 vssd1 vccd1 vccd1 hold5272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5283 _11752_/Y vssd1 vssd1 vccd1 vccd1 _17074_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5294 _16715_/Q vssd1 vssd1 vccd1 vccd1 hold5294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4560 _13645_/X vssd1 vssd1 vccd1 vccd1 _17668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4571 _16701_/Q vssd1 vssd1 vccd1 vccd1 hold4571/X sky130_fd_sc_hd__dlygate4sd3_1
X_10163_ hold1909/X hold3642/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__mux2_1
Xhold4582 _10534_/X vssd1 vssd1 vccd1 vccd1 _16668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4593 _17207_/Q vssd1 vssd1 vccd1 vccd1 hold4593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3870 _12349_/Y vssd1 vssd1 vccd1 vccd1 _17273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3881 _12312_/Y vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14971_ hold1255/X _15006_/B _14970_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _14971_/X
+ sky130_fd_sc_hd__o211a_1
X_10094_ hold1813/X hold3673/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__mux2_1
Xhold3892 _16775_/Q vssd1 vssd1 vccd1 vccd1 hold3892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16710_ _18072_/CLK _16710_/D vssd1 vssd1 vccd1 vccd1 _16710_/Q sky130_fd_sc_hd__dfxtp_1
X_13922_ hold735/X _17769_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 hold736/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17690_ _17722_/CLK _17690_/D vssd1 vssd1 vccd1 vccd1 _17690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _18231_/CLK _16641_/D vssd1 vssd1 vccd1 vccd1 _16641_/Q sky130_fd_sc_hd__dfxtp_1
X_13853_ _17738_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13853_/X sky130_fd_sc_hd__and3_1
X_12804_ _12804_/A _12804_/B vssd1 vssd1 vccd1 vccd1 _17444_/D sky130_fd_sc_hd__and2_1
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16572_ _18206_/CLK _16572_/D vssd1 vssd1 vccd1 vccd1 _16572_/Q sky130_fd_sc_hd__dfxtp_1
X_13784_ hold2091/X hold5102/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__mux2_1
X_10996_ hold5691/X _11789_/B _10995_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10996_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18311_ _18422_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 hold980/A sky130_fd_sc_hd__dfxtp_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ hold949/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__or2_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12756_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _17421_/D sky130_fd_sc_hd__and2_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18243_/CLK hold957/X vssd1 vssd1 vccd1 vccd1 hold956/A sky130_fd_sc_hd__dfxtp_1
X_15454_ _15454_/A _15454_/B vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__and2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _17398_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ hold3351/X _11617_/A2 _11616_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11617_/X
+ sky130_fd_sc_hd__o211a_1
X_14405_ _15193_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18173_ _18205_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15385_ _15385_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__or2_1
X_12597_ _15506_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _17375_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17124_ _18426_/CLK _17124_/D vssd1 vssd1 vccd1 vccd1 _17124_/Q sky130_fd_sc_hd__dfxtp_1
X_11548_ hold4269/X _11735_/B _11547_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14336_ _15231_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 hold519/A vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17055_ _18032_/CLK _17055_/D vssd1 vssd1 vccd1 vccd1 _17055_/Q sky130_fd_sc_hd__dfxtp_1
X_14267_ hold932/X _14266_/B _14266_/Y _15056_/A vssd1 vssd1 vccd1 vccd1 hold933/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ hold5729/X _11765_/B _11478_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11479_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _18413_/CLK _16006_/D vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__dfxtp_1
X_13218_ _17578_/Q _17112_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _15217_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__nand2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13148_/X hold3693/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__mux2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _15855_/Q vssd1 vssd1 vccd1 vccd1 hold1208/X sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ _18063_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1219 _08206_/X vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ _18073_/CLK _16908_/D vssd1 vssd1 vccd1 vccd1 _16908_/Q sky130_fd_sc_hd__dfxtp_1
X_08690_ _12430_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _15966_/D sky130_fd_sc_hd__and2_1
X_17888_ _18427_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_1
X_16839_ _17981_/CLK _16839_/D vssd1 vssd1 vccd1 vccd1 _16839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17503_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09311_ _15099_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09242_ _12777_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _16232_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09173_ hold2590/X _09177_/A2 _09172_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08124_ _15529_/A hold1913/X hold196/X vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08055_ hold2646/X _08082_/B _08054_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _08055_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3100 _17503_/Q vssd1 vssd1 vccd1 vccd1 hold3100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3111 _17504_/Q vssd1 vssd1 vccd1 vccd1 hold3111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3122 _17430_/Q vssd1 vssd1 vccd1 vccd1 hold3122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3133 _10605_/Y vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3144 _16523_/Q vssd1 vssd1 vccd1 vccd1 hold3144/X sky130_fd_sc_hd__clkbuf_2
Xhold2410 _14729_/X vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3155 _12352_/Y vssd1 vssd1 vccd1 vccd1 _17274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3166 _12294_/Y vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2421 _17881_/Q vssd1 vssd1 vccd1 vccd1 hold2421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 _08396_/X vssd1 vssd1 vccd1 vccd1 _15828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3177 _16361_/Q vssd1 vssd1 vccd1 vccd1 hold3177/X sky130_fd_sc_hd__dlygate4sd3_1
X_08957_ hold136/X hold304/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__mux2_1
Xhold3188 _16520_/Q vssd1 vssd1 vccd1 vccd1 hold3188/X sky130_fd_sc_hd__buf_2
Xhold2443 _18441_/Q vssd1 vssd1 vccd1 vccd1 hold2443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2454 _14657_/X vssd1 vssd1 vccd1 vccd1 _18121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3199 _17461_/Q vssd1 vssd1 vccd1 vccd1 hold3199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1720 _18172_/Q vssd1 vssd1 vccd1 vccd1 hold1720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2465 _08332_/X vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1731 _13039_/X vssd1 vssd1 vccd1 vccd1 _17523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2476 _18113_/Q vssd1 vssd1 vccd1 vccd1 hold2476/X sky130_fd_sc_hd__dlygate4sd3_1
X_07908_ _14866_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__or2_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2487 _18279_/Q vssd1 vssd1 vccd1 vccd1 hold2487/X sky130_fd_sc_hd__dlygate4sd3_1
X_08888_ hold443/X hold564/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__mux2_1
Xhold1742 _16189_/Q vssd1 vssd1 vccd1 vccd1 hold1742/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2498 _14919_/X vssd1 vssd1 vccd1 vccd1 _18246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1753 _09095_/X vssd1 vssd1 vccd1 vccd1 _16162_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1764 _15156_/X vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1775 hold5823/X vssd1 vssd1 vccd1 vccd1 _13030_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _14511_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__or2_1
Xhold1786 _15882_/Q vssd1 vssd1 vccd1 vccd1 hold1786/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1797 _18091_/Q vssd1 vssd1 vccd1 vccd1 hold1797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10850_ hold1118/X hold4341/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _18240_/Q _13086_/A _09998_/C vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ hold2578/X hold4131/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10782_/B sky130_fd_sc_hd__mux2_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ hold1874/X _17351_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__mux2_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ hold78/X _12509_/A2 _12505_/A3 _12450_/X _12420_/A vssd1 vssd1 vccd1 vccd1
+ hold79/A sky130_fd_sc_hd__o311a_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11402_ hold2026/X _16958_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _11403_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ hold2078/X hold609/X _15169_/X _15482_/A vssd1 vssd1 vccd1 vccd1 _15170_/X
+ sky130_fd_sc_hd__o211a_1
X_12382_ _15244_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _17284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_90 hold5876/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ hold2666/X hold587/X _14120_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ hold2895/X hold3382/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14052_ _14786_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11264_ hold2276/X hold3790/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11265_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5080 _16787_/Q vssd1 vssd1 vccd1 vccd1 hold5080/X sky130_fd_sc_hd__dlygate4sd3_1
X_13003_ _14897_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__nor2_2
X_10215_ _10548_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__or2_1
Xhold5091 _11686_/X vssd1 vssd1 vccd1 vccd1 _17052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_11195_ _16889_/Q _11762_/B _11762_/C vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4390 _11896_/X vssd1 vssd1 vccd1 vccd1 _17122_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17811_ _17893_/CLK hold994/X vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__dfxtp_1
X_10146_ _10485_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17742_ _17742_/CLK _17742_/D vssd1 vssd1 vccd1 vccd1 _17742_/Q sky130_fd_sc_hd__dfxtp_1
X_14954_ hold730/X _14962_/B vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__or2_1
X_10077_ _10563_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10077_/X sky130_fd_sc_hd__or2_1
X_13905_ _13905_/A _13905_/B vssd1 vssd1 vccd1 vccd1 _17760_/D sky130_fd_sc_hd__and2_1
X_17673_ _17737_/CLK _17673_/D vssd1 vssd1 vccd1 vccd1 _17673_/Q sky130_fd_sc_hd__dfxtp_1
X_14885_ hold758/X _14882_/B _14884_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 hold759/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16624_ _18206_/CLK _16624_/D vssd1 vssd1 vccd1 vccd1 _16624_/Q sky130_fd_sc_hd__dfxtp_1
X_13836_ hold3894/X _13776_/A _13835_/X vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16555_ _18392_/CLK _16555_/D vssd1 vssd1 vccd1 vccd1 _16555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ hold2921/X _16817_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15506_ _15506_/A _15506_/B vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__and2_1
X_12718_ hold2455/X _17417_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _18339_/CLK _16486_/D vssd1 vssd1 vccd1 vccd1 _16486_/Q sky130_fd_sc_hd__dfxtp_1
X_13698_ _13767_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__or2_1
X_18225_ _18225_/CLK hold819/X vssd1 vssd1 vccd1 vccd1 hold818/A sky130_fd_sc_hd__dfxtp_1
X_15437_ hold304/X _09392_/B _09392_/C hold321/X vssd1 vssd1 vccd1 vccd1 _15437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ hold2407/X _17394_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _18216_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
X_15368_ hold649/X _15484_/A2 _15451_/A2 hold663/X vssd1 vssd1 vccd1 vccd1 _15368_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ _17865_/CLK _17107_/D vssd1 vssd1 vccd1 vccd1 _17107_/Q sky130_fd_sc_hd__dfxtp_1
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319_ hold1553/X _14326_/B _14318_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14319_/X
+ sky130_fd_sc_hd__o211a_1
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _18268_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15299_ hold702/X _15485_/A2 _15447_/B1 hold680/X _15298_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _18051_/CLK _17038_/D vssd1 vssd1 vccd1 vccd1 _17038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout807 _15208_/C1 vssd1 vssd1 vccd1 vccd1 _15216_/C1 sky130_fd_sc_hd__buf_4
X_09860_ hold1246/X _16444_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14392_/A sky130_fd_sc_hd__buf_4
Xfanout829 _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/C1 sky130_fd_sc_hd__buf_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _09003_/A _08811_/B vssd1 vssd1 vccd1 vccd1 _16024_/D sky130_fd_sc_hd__and2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ hold2856/X _16421_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _15216_/X vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _17918_/Q vssd1 vssd1 vccd1 vccd1 hold1016/X sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _12422_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _15991_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _15783_/Q vssd1 vssd1 vccd1 vccd1 hold1027/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 hold128/X vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _15676_/Q vssd1 vssd1 vccd1 vccd1 hold1049/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ hold32/X hold330/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ hold2384/X _09216_/B _09224_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _09225_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_256_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17732_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09156_ _15105_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08107_ _08161_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _15692_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09087_ hold2858/X _09119_/A2 _09086_/X _12987_/A vssd1 vssd1 vccd1 vccd1 _09087_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ hold1405/X _08033_/B _08037_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _08038_/X
+ sky130_fd_sc_hd__o211a_1
Xhold850 hold850/A vssd1 vssd1 vccd1 vccd1 input54/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 hold861/A vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold872 hold872/A vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__clkbuf_16
Xhold894 hold894/A vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _11155_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10000_/Y sky130_fd_sc_hd__nor2_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _09989_/A _09998_/B _09998_/C vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__and3_1
Xhold2240 _08034_/X vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 _09101_/X vssd1 vssd1 vccd1 vccd1 _16165_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2262 _18306_/Q vssd1 vssd1 vccd1 vccd1 hold2262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2273 _14989_/X vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2284 _14865_/X vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1550 _17521_/Q vssd1 vssd1 vccd1 vccd1 hold1550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2295 _15653_/Q vssd1 vssd1 vccd1 vccd1 hold2295/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1561 _17785_/Q vssd1 vssd1 vccd1 vccd1 hold1561/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1572 _14929_/X vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11951_ hold2336/X hold4765/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1583 _14887_/X vssd1 vssd1 vccd1 vccd1 _18232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 _14857_/X vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _11121_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__or2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _15225_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__or2_1
X_11882_ _15710_/Q hold3731/X _13871_/C vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__mux2_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13621_ hold4959/X _13805_/B _13620_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__o211a_1
X_10833_ _11121_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10833_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16340_ _18363_/CLK _16340_/D vssd1 vssd1 vccd1 vccd1 _16340_/Q sky130_fd_sc_hd__dfxtp_1
X_13552_ hold4838/X _13856_/B _13551_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13552_/X
+ sky130_fd_sc_hd__o211a_1
X_10764_ _11136_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12503_ hold29/X _08598_/B _08999_/B _12502_/X _09047_/A vssd1 vssd1 vccd1 vccd1
+ hold30/A sky130_fd_sc_hd__o311a_1
XFILLER_0_165_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13483_ hold4633/X _13832_/B _13482_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13483_/X
+ sky130_fd_sc_hd__o211a_1
X_16271_ _17375_/CLK _16271_/D vssd1 vssd1 vccd1 vccd1 _16271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10695_ _11115_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ _18431_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ hold930/X _15221_/B _15221_/Y _15024_/A vssd1 vssd1 vccd1 vccd1 hold931/A
+ sky130_fd_sc_hd__o211a_1
X_12434_ _15374_/A _12434_/B vssd1 vssd1 vccd1 vccd1 _17310_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _15207_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12365_ _17279_/Q _12374_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12365_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11316_ _12246_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__or2_1
X_14104_ _15123_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__or2_1
X_15084_ hold1587/X _15113_/B _15083_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _15084_/X
+ sky130_fd_sc_hd__o211a_1
X_12296_ _17256_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__and3_1
X_14035_ hold1939/X _14040_/B _14034_/Y _13909_/A vssd1 vssd1 vccd1 vccd1 _14035_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11247_ _11631_/A _11247_/B vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11178_ hold3648/X _11082_/A _11177_/X vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__a21oi_1
X_10129_ hold4083/X _10631_/B _10128_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15986_ _17525_/CLK _15986_/D vssd1 vssd1 vccd1 vccd1 hold631/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17725_/CLK _17725_/D vssd1 vssd1 vccd1 vccd1 _17725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14937_ hold2787/X _14952_/B _14936_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14937_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17656_ _17725_/CLK _17656_/D vssd1 vssd1 vccd1 vccd1 _17656_/Q sky130_fd_sc_hd__dfxtp_1
X_14868_ _15099_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__or2_1
X_16607_ _18131_/CLK _16607_/D vssd1 vssd1 vccd1 vccd1 _16607_/Q sky130_fd_sc_hd__dfxtp_1
X_13819_ _13822_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _13819_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_5_24__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_24__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17587_ _17747_/CLK _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ hold1330/X _14822_/B _14798_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14799_/X
+ sky130_fd_sc_hd__o211a_1
X_16538_ _18224_/CLK _16538_/D vssd1 vssd1 vccd1 vccd1 _16538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ _18382_/CLK _16469_/D vssd1 vssd1 vccd1 vccd1 _16469_/Q sky130_fd_sc_hd__dfxtp_1
X_09010_ hold41/X hold388/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ _18208_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5805 output74/X vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_12
X_18139_ _18395_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5816 _18406_/Q vssd1 vssd1 vccd1 vccd1 hold5816/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5827 hold5937/X vssd1 vssd1 vccd1 vccd1 hold5827/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5838 _16280_/Q vssd1 vssd1 vccd1 vccd1 hold5838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold262/X vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5849 hold5849/A vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_12
Xhold135 input7/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 data_in[23] vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold46/X vssd1 vssd1 vccd1 vccd1 input34/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09912_ _09924_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__or2_1
Xhold179 hold11/X vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__buf_4
XFILLER_0_10_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout604 _15484_/B1 vssd1 vssd1 vccd1 vccd1 _09386_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout615 _09358_/Y vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__clkbuf_8
Xfanout626 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15490_/A1 sky130_fd_sc_hd__buf_6
X_09843_ _09987_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__or2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout637 _12849_/A vssd1 vssd1 vccd1 vccd1 _12789_/A sky130_fd_sc_hd__buf_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout648 _12885_/A vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__buf_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout659 fanout660/X vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__clkbuf_4
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _10506_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__or2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ hold14/X hold200/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _15454_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _15950_/D sky130_fd_sc_hd__and2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08887_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _15917_/D sky130_fd_sc_hd__and2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09208_ _15537_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _10574_/A _11177_/B _10479_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10480_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09139_ hold2586/X _09177_/A2 _09138_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12150_ _12282_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ hold5389/X _11753_/B _11100_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11101_/X
+ sky130_fd_sc_hd__o211a_1
X_12081_ _12279_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 hold680/A vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold691 hold691/A vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ hold5662/X _11789_/B _11031_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _11032_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _17669_/CLK _15840_/D vssd1 vssd1 vccd1 vccd1 _15840_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _18149_/Q vssd1 vssd1 vccd1 vccd1 hold2070/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2081 _14275_/X vssd1 vssd1 vccd1 vccd1 _17938_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 _08216_/X vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _17722_/CLK _15771_/D vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ hold3111/X _12982_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12983_/X sky130_fd_sc_hd__mux2_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1380 _14917_/X vssd1 vssd1 vccd1 vccd1 _18245_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17510_ _17511_/CLK _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _15169_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14722_/X sky130_fd_sc_hd__or2_1
Xhold1391 _18363_/Q vssd1 vssd1 vccd1 vccd1 hold1391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _12267_/A _11934_/B vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17448_/CLK _17441_/D vssd1 vssd1 vccd1 vccd1 _17441_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_178_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18190_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14653_ hold2203/X _14664_/B _14652_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14653_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ _13749_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__or2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ hold2201/X hold4117/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18243_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17372_ _18431_/CLK _17372_/D vssd1 vssd1 vccd1 vccd1 _17372_/Q sky130_fd_sc_hd__dfxtp_1
X_10816_ hold5687/X _11789_/B _10815_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _10816_/X
+ sky130_fd_sc_hd__o211a_1
X_11796_ hold3952/X _12246_/A _11795_/X vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__a21oi_1
X_14584_ _15193_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16323_ _17503_/CLK _16323_/D vssd1 vssd1 vccd1 vccd1 _16323_/Q sky130_fd_sc_hd__dfxtp_1
X_13535_ hold913/X hold3357/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ hold5329/X _11765_/B _10746_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _10747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ _17487_/CLK _16254_/D vssd1 vssd1 vccd1 vccd1 _16254_/Q sky130_fd_sc_hd__dfxtp_1
X_13466_ hold845/X _17609_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13467_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ hold5586/X _11156_/B _10677_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10678_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _15205_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__or2_1
X_12417_ hold219/X _17302_/Q _12443_/S vssd1 vssd1 vccd1 vccd1 hold547/A sky130_fd_sc_hd__mux2_1
X_16185_ _18451_/CLK _16185_/D vssd1 vssd1 vccd1 vccd1 _16185_/Q sky130_fd_sc_hd__dfxtp_1
X_13397_ hold1240/X hold3931/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15136_ hold2965/X hold609/X _15135_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15136_/X
+ sky130_fd_sc_hd__o211a_1
X_12348_ hold3868/X _12255_/A _12347_/X vssd1 vssd1 vccd1 vccd1 _12348_/Y sky130_fd_sc_hd__a21oi_1
X_12279_ _12279_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__or2_1
X_15067_ _15229_/A hold2090/X hold302/X vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_5_8__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_8__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_14018_ _15525_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15969_ _17522_/CLK _15969_/D vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_1
X_08510_ hold1786/X _08503_/Y _08509_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08510_/X
+ sky130_fd_sc_hd__o211a_1
X_17708_ _17708_/CLK _17708_/D vssd1 vssd1 vccd1 vccd1 _17708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ _13030_/A _13043_/C _17518_/Q vssd1 vssd1 vccd1 vccd1 _13055_/C sky130_fd_sc_hd__and3_4
X_08441_ _14728_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__or2_1
X_17639_ _17735_/CLK _17639_/D vssd1 vssd1 vccd1 vccd1 _17639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ hold265/A _15818_/Q hold122/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__mux2_1
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5602 _16360_/Q vssd1 vssd1 vccd1 vccd1 hold5602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5613 _09703_/X vssd1 vssd1 vccd1 vccd1 _16391_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5624 _11041_/X vssd1 vssd1 vccd1 vccd1 _16837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5635 _16400_/Q vssd1 vssd1 vccd1 vccd1 hold5635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4901 _16647_/Q vssd1 vssd1 vccd1 vccd1 hold4901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5646 _11092_/X vssd1 vssd1 vccd1 vccd1 _16854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4912 _11338_/X vssd1 vssd1 vccd1 vccd1 _16936_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5657 _16792_/Q vssd1 vssd1 vccd1 vccd1 hold5657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4923 _17271_/Q vssd1 vssd1 vccd1 vccd1 hold4923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5668 _16831_/Q vssd1 vssd1 vccd1 vccd1 hold5668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4934 _12250_/X vssd1 vssd1 vccd1 vccd1 _17240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5679 _16783_/Q vssd1 vssd1 vccd1 vccd1 hold5679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4945 _17186_/Q vssd1 vssd1 vccd1 vccd1 hold4945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4956 _13390_/X vssd1 vssd1 vccd1 vccd1 _17583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4967 _17059_/Q vssd1 vssd1 vccd1 vccd1 hold4967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4978 _10378_/X vssd1 vssd1 vccd1 vccd1 _16616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout401 _14411_/B vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__clkbuf_8
Xfanout412 _14206_/B vssd1 vssd1 vccd1 vccd1 _14214_/B sky130_fd_sc_hd__clkbuf_8
Xhold4989 _17558_/Q vssd1 vssd1 vccd1 vccd1 hold4989/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout423 _14000_/Y vssd1 vssd1 vccd1 vccd1 _14036_/B sky130_fd_sc_hd__buf_6
Xfanout434 _13052_/X vssd1 vssd1 vccd1 vccd1 _13311_/A1 sky130_fd_sc_hd__buf_8
Xfanout445 _12353_/C vssd1 vssd1 vccd1 vccd1 _12356_/C sky130_fd_sc_hd__clkbuf_8
Xfanout456 _11171_/C vssd1 vssd1 vccd1 vccd1 _11747_/C sky130_fd_sc_hd__clkbuf_8
Xfanout467 fanout484/X vssd1 vssd1 vccd1 vccd1 _13886_/C sky130_fd_sc_hd__clkbuf_8
X_09826_ hold5610/X _11201_/B _09825_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _09826_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout478 _11672_/S vssd1 vssd1 vccd1 vccd1 _12341_/C sky130_fd_sc_hd__clkbuf_8
Xfanout489 _10874_/S vssd1 vssd1 vccd1 vccd1 _09998_/C sky130_fd_sc_hd__clkbuf_8
X_09757_ hold5359/X _10025_/B _09756_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09757_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _12402_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _15975_/D sky130_fd_sc_hd__and2_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ hold4688/X _10070_/B _09687_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09688_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_271_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17865_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ hold5/X hold217/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__mux2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_200_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18060_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_166_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11744_/A _11741_/B _11649_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11650_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10601_ _16691_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__and3_1
XFILLER_0_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ hold5381/X _12338_/B _11580_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11581_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ hold1304/X hold4449/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__mux2_1
X_13320_ _13713_/A _13320_/B vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10463_ hold2875/X _16645_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__mux2_1
X_13251_ _13250_/X _16924_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ hold4551/X _13811_/B _12201_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _12202_/X
+ sky130_fd_sc_hd__o211a_1
X_13182_ _13182_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__or2_1
X_10394_ hold1495/X _16622_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__mux2_1
X_12133_ hold4781/X _12314_/B _12132_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12133_/X
+ sky130_fd_sc_hd__o211a_1
X_17990_ _18054_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12064_ hold5030/X _12347_/B _12063_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12064_/X
+ sky130_fd_sc_hd__o211a_1
X_16941_ _17856_/CLK _16941_/D vssd1 vssd1 vccd1 vccd1 _16941_/Q sky130_fd_sc_hd__dfxtp_1
X_11015_ hold820/X hold4405/X _11219_/C vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__mux2_1
X_16872_ _18043_/CLK _16872_/D vssd1 vssd1 vccd1 vccd1 _16872_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _17734_/CLK _15823_/D vssd1 vssd1 vccd1 vccd1 _15823_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _17715_/CLK _15754_/D vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _12984_/A _12966_/B vssd1 vssd1 vccd1 vccd1 _17498_/D sky130_fd_sc_hd__and2_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ hold2938/X _14720_/B _14704_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ hold4971/X _12299_/B _11916_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__o211a_1
X_15685_ _17583_/CLK _15685_/D vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _15506_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _17475_/D sky130_fd_sc_hd__and2_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17424_ _17629_/CLK _17424_/D vssd1 vssd1 vccd1 vccd1 _17424_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _15191_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14636_/X sky130_fd_sc_hd__or2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ hold3427/X _13871_/B _11847_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _11848_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17516_/CLK _17355_/D vssd1 vssd1 vccd1 vccd1 _17355_/Q sky130_fd_sc_hd__dfxtp_1
X_14567_ _15191_/A _14557_/Y hold935/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 hold936/A
+ sky130_fd_sc_hd__o211a_1
X_11779_ _12301_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _17511_/CLK _16306_/D vssd1 vssd1 vccd1 vccd1 _16306_/Q sky130_fd_sc_hd__dfxtp_1
X_13518_ _13710_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17286_ _18409_/CLK _17286_/D vssd1 vssd1 vccd1 vccd1 _17286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ hold2967/X _14487_/B _14497_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _14498_/X
+ sky130_fd_sc_hd__o211a_1
X_16237_ _17419_/CLK _16237_/D vssd1 vssd1 vccd1 vccd1 _16237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13449_ _13737_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17522_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4208 _13726_/X vssd1 vssd1 vccd1 vccd1 _17695_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16168_ _17506_/CLK hold763/X vssd1 vssd1 vccd1 vccd1 hold762/A sky130_fd_sc_hd__dfxtp_1
Xhold4219 _11920_/X vssd1 vssd1 vccd1 vccd1 _17130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15119_ _15227_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15119_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3507 _17172_/Q vssd1 vssd1 vccd1 vccd1 hold3507/X sky130_fd_sc_hd__dlygate4sd3_1
X_08990_ _09047_/A _08990_/B vssd1 vssd1 vccd1 vccd1 _16112_/D sky130_fd_sc_hd__and2_1
X_16099_ _17531_/CLK _16099_/D vssd1 vssd1 vccd1 vccd1 _16099_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3518 _12809_/X vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3529 _16511_/Q vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07941_ hold1484/X _07991_/A2 _07940_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07941_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2806 _08063_/X vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2817 _15098_/X vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 _18054_/Q vssd1 vssd1 vccd1 vccd1 hold2828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2839 _14981_/X vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07872_ hold1960/X _07869_/B _07871_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07872_/X
+ sky130_fd_sc_hd__o211a_1
X_09611_ _18274_/Q hold3177/X _09998_/C vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09542_ hold1571/X _13174_/A _10022_/C vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09473_ _09477_/C _09481_/B _09473_/C vssd1 vssd1 vccd1 vccd1 _16318_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08424_ hold833/X _08433_/B _08423_/X _08381_/A vssd1 vssd1 vccd1 vccd1 hold834/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _15809_/D sky130_fd_sc_hd__and2_1
XFILLER_0_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08286_ hold1242/X _08336_/A2 _08285_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08286_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5410 _11374_/X vssd1 vssd1 vccd1 vccd1 _16948_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5421 _16818_/Q vssd1 vssd1 vccd1 vccd1 hold5421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5432 _11089_/X vssd1 vssd1 vccd1 vccd1 _16853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5443 _16953_/Q vssd1 vssd1 vccd1 vccd1 hold5443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5454 _16396_/Q vssd1 vssd1 vccd1 vccd1 hold5454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4720 _17698_/Q vssd1 vssd1 vccd1 vccd1 hold4720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5465 _11116_/X vssd1 vssd1 vccd1 vccd1 _16862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5476 _16421_/Q vssd1 vssd1 vccd1 vccd1 hold5476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4731 _17712_/Q vssd1 vssd1 vccd1 vccd1 hold4731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4742 _15373_/X vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5487 _11404_/X vssd1 vssd1 vccd1 vccd1 _16958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4753 _16482_/Q vssd1 vssd1 vccd1 vccd1 hold4753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5498 _16371_/Q vssd1 vssd1 vccd1 vccd1 hold5498/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4764 _11899_/X vssd1 vssd1 vccd1 vccd1 _17123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4775 _17689_/Q vssd1 vssd1 vccd1 vccd1 hold4775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4786 _12127_/X vssd1 vssd1 vccd1 vccd1 _17199_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 _10001_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__buf_4
Xhold4797 _17188_/Q vssd1 vssd1 vccd1 vccd1 hold4797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout231 _10610_/B vssd1 vssd1 vccd1 vccd1 _10643_/B sky130_fd_sc_hd__buf_4
XFILLER_0_79_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout242 _10649_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__clkbuf_8
Xfanout253 _12210_/A vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__buf_4
Xfanout264 _11616_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__clkbuf_4
Xfanout275 _13770_/A vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__buf_2
Xfanout286 _11688_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__clkbuf_4
X_09809_ hold2258/X _16427_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__mux2_1
Xfanout297 fanout298/X vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__buf_4
X_12820_ hold1830/X hold3083/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12751_ hold1863/X _17428_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__mux2_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ hold1533/X _17058_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__mux2_1
X_15470_ _16051_/Q _09392_/C _15467_/X vssd1 vssd1 vccd1 vccd1 _15471_/D sky130_fd_sc_hd__a21o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ hold2734/X _17405_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _15535_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__or2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11633_ hold2834/X _17035_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _17274_/CLK _17140_/D vssd1 vssd1 vccd1 vccd1 _17140_/Q sky130_fd_sc_hd__dfxtp_1
X_14352_ _14352_/A hold827/X vssd1 vssd1 vccd1 vccd1 hold828/A sky130_fd_sc_hd__and2_1
XFILLER_0_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ hold983/X _17012_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ _13311_/A1 _13301_/X _13302_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__or2_1
X_17071_ _17887_/CLK _17071_/D vssd1 vssd1 vccd1 vccd1 _17071_/Q sky130_fd_sc_hd__dfxtp_1
X_11495_ hold991/X _16989_/Q _12338_/C vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__mux2_1
X_14283_ hold2915/X _14272_/B _14282_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14283_/X
+ sky130_fd_sc_hd__o211a_1
X_16022_ _17323_/CLK _16022_/D vssd1 vssd1 vccd1 vccd1 hold644/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ _10542_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__or2_1
X_13234_ _17580_/Q _17114_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13164_/X hold5899/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__mux2_1
X_10377_ _10491_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__or2_1
X_12116_ hold1861/X _17196_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__mux2_1
X_13096_ _13089_/X _13095_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17530_/D sky130_fd_sc_hd__o21a_1
X_17973_ _18032_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12047_ hold1983/X _17173_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _12048_/B sky130_fd_sc_hd__mux2_1
X_16924_ _17890_/CLK _16924_/D vssd1 vssd1 vccd1 vccd1 _16924_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_193_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16855_ _18067_/CLK _16855_/D vssd1 vssd1 vccd1 vccd1 _16855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15806_ _17745_/CLK _15806_/D vssd1 vssd1 vccd1 vccd1 hold977/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_122_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ _18053_/CLK _16786_/D vssd1 vssd1 vccd1 vccd1 _16786_/Q sky130_fd_sc_hd__dfxtp_1
X_13998_ _14786_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _17708_/CLK _15737_/D vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfxtp_1
X_12949_ hold2752/X hold3583/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__mux2_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _18456_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
X_15668_ _17128_/CLK _15668_/D vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17407_ _18458_/CLK _17407_/D vssd1 vssd1 vccd1 vccd1 _17407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14619_ hold1909/X _14612_/B _14618_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14619_/X
+ sky130_fd_sc_hd__o211a_1
X_18387_ _18395_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _17282_/CLK _15599_/D vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ hold335/X hold516/X hold196/X vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__mux2_1
X_17338_ _17341_/CLK hold141/X vssd1 vssd1 vccd1 vccd1 _17338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ hold2040/X _08082_/B _08070_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _08071_/X
+ sky130_fd_sc_hd__o211a_1
X_17269_ _17777_/CLK _17269_/D vssd1 vssd1 vccd1 vccd1 _17269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4005 _10630_/Y vssd1 vssd1 vccd1 vccd1 _16700_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4016 _16641_/Q vssd1 vssd1 vccd1 vccd1 hold4016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4027 _11047_/X vssd1 vssd1 vccd1 vccd1 _16839_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4038 _15293_/X vssd1 vssd1 vccd1 vccd1 _15294_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4049 _17688_/Q vssd1 vssd1 vccd1 vccd1 hold4049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3304 _12857_/X vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3315 _17152_/Q vssd1 vssd1 vccd1 vccd1 hold3315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3326 _16604_/Q vssd1 vssd1 vccd1 vccd1 hold3326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3337 _13345_/X vssd1 vssd1 vccd1 vccd1 _17568_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08973_ hold17/X hold84/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__mux2_1
Xhold2603 _18208_/Q vssd1 vssd1 vccd1 vccd1 hold2603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3348 _11986_/X vssd1 vssd1 vccd1 vccd1 _17152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3359 _09961_/X vssd1 vssd1 vccd1 vccd1 _16477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2614 _18022_/Q vssd1 vssd1 vccd1 vccd1 hold2614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold75/X vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__buf_4
Xhold2625 _09193_/X vssd1 vssd1 vccd1 vccd1 _16208_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _15547_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07924_/Y sky130_fd_sc_hd__nand2_1
Xhold2636 _09089_/X vssd1 vssd1 vccd1 vccd1 _16159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1902 _08028_/X vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 _08055_/X vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _15701_/Q vssd1 vssd1 vccd1 vccd1 hold1913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _17813_/Q vssd1 vssd1 vccd1 vccd1 hold2658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 _09163_/X vssd1 vssd1 vccd1 vccd1 _16194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 _14771_/X vssd1 vssd1 vccd1 vccd1 _18176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 _08326_/X vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _15533_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__or2_1
Xhold1946 _09213_/X vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 _14219_/X vssd1 vssd1 vccd1 vccd1 _17911_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _15688_/Q vssd1 vssd1 vccd1 vccd1 hold1968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1979 _17913_/Q vssd1 vssd1 vccd1 vccd1 hold1979/X sky130_fd_sc_hd__dlygate4sd3_1
X_07786_ _16287_/Q vssd1 vssd1 vccd1 vccd1 _07786_/Y sky130_fd_sc_hd__inv_2
X_09525_ _09933_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09463_/D
+ sky130_fd_sc_hd__and4_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _15521_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09387_ _15471_/A _09386_/X _18460_/Q vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ hold606/A hold298/A _09399_/C vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__or3_1
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08269_ hold1807/X _08268_/B _08268_/Y _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08269_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ hold4271/X _10589_/B _10299_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11280_ _11670_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11280_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5240 _12330_/Y vssd1 vssd1 vccd1 vccd1 _12331_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10231_ hold3219/X _10637_/B _10230_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5251 _16725_/Q vssd1 vssd1 vccd1 vccd1 hold5251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5262 _11206_/Y vssd1 vssd1 vccd1 vccd1 _16892_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5273 _11787_/Y vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5284 _16329_/Q vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4550 _09859_/X vssd1 vssd1 vccd1 vccd1 _16443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5295 _11154_/Y vssd1 vssd1 vccd1 vccd1 _11155_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4561 _16633_/Q vssd1 vssd1 vccd1 vccd1 hold4561/X sky130_fd_sc_hd__dlygate4sd3_1
X_10162_ hold4359/X _10640_/B _10161_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10162_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4572 _10537_/X vssd1 vssd1 vccd1 vccd1 _16669_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4583 _17090_/Q vssd1 vssd1 vccd1 vccd1 hold4583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4594 _12055_/X vssd1 vssd1 vccd1 vccd1 _17175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3860 _09529_/X vssd1 vssd1 vccd1 vccd1 _16333_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3871 _16931_/Q vssd1 vssd1 vccd1 vccd1 hold3871/X sky130_fd_sc_hd__dlygate4sd3_1
X_14970_ _14970_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__or2_1
X_10093_ hold4093/X _10571_/B _10092_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _10093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3882 _12313_/Y vssd1 vssd1 vccd1 vccd1 _17261_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3893 _10759_/X vssd1 vssd1 vccd1 vccd1 _16743_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13921_ _13935_/A _13921_/B vssd1 vssd1 vccd1 vccd1 _17768_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16640_ _18198_/CLK _16640_/D vssd1 vssd1 vccd1 vccd1 _16640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _13888_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__nor2_1
X_12803_ hold3523/X _12802_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12804_/B sky130_fd_sc_hd__mux2_1
X_16571_ _18225_/CLK _16571_/D vssd1 vssd1 vccd1 vccd1 _16571_/Q sky130_fd_sc_hd__dfxtp_1
X_13783_ hold5052/X _13880_/B _13782_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13783_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10995_ _11694_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10995_/X sky130_fd_sc_hd__or2_1
X_18310_ _18420_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ hold2481/X _15560_/A2 _15521_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _15522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ hold3085/X _12733_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12735_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/CLK hold658/X vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ _15490_/A1 _15445_/X _15452_/X _15490_/B1 _18421_/Q vssd1 vssd1 vccd1 vccd1
+ _15453_/X sky130_fd_sc_hd__a32o_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12665_ hold3055/X _12664_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__mux2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ hold1546/X hold209/X _14403_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14404_/X
+ sky130_fd_sc_hd__o211a_1
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__or2_1
X_18172_ _18228_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
X_15384_ _15482_/A _15384_/B vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__and2_1
XFILLER_0_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12596_ hold3375/X _12595_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17123_ _17281_/CLK _17123_/D vssd1 vssd1 vccd1 vccd1 _17123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ hold2427/X _14326_/B _14334_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _14335_/X
+ sky130_fd_sc_hd__o211a_1
X_11547_ _11640_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold509 hold509/A vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ _17870_/CLK _17054_/D vssd1 vssd1 vccd1 vccd1 _17054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _15215_/A _14266_/B vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__nand2_1
X_11478_ _11670_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ _18416_/CLK _16005_/D vssd1 vssd1 vccd1 vccd1 _16005_/Q sky130_fd_sc_hd__dfxtp_1
X_13217_ _13217_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10429_ hold4665/X _10637_/B _10428_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10429_/X
+ sky130_fd_sc_hd__o211a_1
X_14197_ hold2050/X _14198_/B _14196_/Y _13931_/A vssd1 vssd1 vccd1 vccd1 _14197_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ hold3604/X _13147_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__mux2_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17634_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _18053_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
X_13079_ _13183_/A1 _13077_/X _13078_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13079_/X
+ sky130_fd_sc_hd__o211a_2
Xhold1209 _08453_/X vssd1 vssd1 vccd1 vccd1 _15855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16907_ _17852_/CLK _16907_/D vssd1 vssd1 vccd1 vccd1 _16907_/Q sky130_fd_sc_hd__dfxtp_1
X_17887_ _17887_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_1
X_16838_ _18009_/CLK _16838_/D vssd1 vssd1 vccd1 vccd1 _16838_/Q sky130_fd_sc_hd__dfxtp_1
X_16769_ _18069_/CLK _16769_/D vssd1 vssd1 vccd1 vccd1 _16769_/Q sky130_fd_sc_hd__dfxtp_1
X_09310_ hold1648/X _09325_/B _09309_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _15517_/A hold997/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__mux2_1
X_18439_ _18454_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_90_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17531_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09172_ hold800/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08123_ _08133_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__and2_1
XFILLER_0_145_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ _15513_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3101 _12980_/X vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3112 _12983_/X vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3123 _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3134 _10606_/Y vssd1 vssd1 vccd1 vccd1 _16692_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 _10578_/Y vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2400 _07842_/X vssd1 vssd1 vccd1 vccd1 _15566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 _15729_/Q vssd1 vssd1 vccd1 vccd1 hold2411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3156 _16911_/Q vssd1 vssd1 vccd1 vccd1 hold3156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 _12295_/Y vssd1 vssd1 vccd1 vccd1 _17255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2422 _14155_/X vssd1 vssd1 vccd1 vccd1 _17881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08956_ _15473_/A hold163/X vssd1 vssd1 vccd1 vccd1 _16095_/D sky130_fd_sc_hd__and2_1
Xhold2433 _18295_/Q vssd1 vssd1 vccd1 vccd1 hold2433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3178 _09517_/X vssd1 vssd1 vccd1 vccd1 _16329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3189 _10569_/Y vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2444 _15526_/X vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1710 _16215_/Q vssd1 vssd1 vccd1 vccd1 hold1710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2455 _16237_/Q vssd1 vssd1 vccd1 vccd1 hold2455/X sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ hold2076/X _07918_/B _07906_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07907_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2466 _16263_/Q vssd1 vssd1 vccd1 vccd1 hold2466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1721 _14763_/X vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2477 _14641_/X vssd1 vssd1 vccd1 vccd1 _18113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1732 _18108_/Q vssd1 vssd1 vccd1 vccd1 hold1732/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _16061_/D sky130_fd_sc_hd__and2_1
Xhold1743 _09153_/X vssd1 vssd1 vccd1 vccd1 _16189_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2488 _14987_/X vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2499 _18130_/Q vssd1 vssd1 vccd1 vccd1 hold2499/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _17820_/Q vssd1 vssd1 vccd1 vccd1 hold1754/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1765 _15737_/Q vssd1 vssd1 vccd1 vccd1 hold1765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1776 _13029_/X vssd1 vssd1 vccd1 vccd1 _13031_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ hold1675/X _07865_/B _07837_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _07838_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1787 _08510_/X vssd1 vssd1 vccd1 vccd1 _15882_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 _14595_/X vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ hold5568/X _09998_/B _09507_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09508_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ hold3983/X _10780_/A2 _10779_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _10780_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ hold1601/X _07804_/A _15334_/A _09438_/X vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _17318_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11401_ hold5456/X _12338_/B _11400_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11401_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12381_ hold23/X hold475/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_80 _15207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_91 hold5901/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14854_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ hold4629/X _12305_/B _11331_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14051_ hold1349/X _14036_/B _14050_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14051_/X
+ sky130_fd_sc_hd__o211a_1
X_11263_ hold4524/X _11741_/B _11262_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5070 _16998_/Q vssd1 vssd1 vccd1 vccd1 hold5070/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5081 _10795_/X vssd1 vssd1 vccd1 vccd1 _16755_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _17510_/D sky130_fd_sc_hd__and2_1
X_10214_ hold1708/X _16562_/Q _10643_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__mux2_1
Xhold5092 _17682_/Q vssd1 vssd1 vccd1 vccd1 hold5092/X sky130_fd_sc_hd__dlygate4sd3_1
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11194_/Y sky130_fd_sc_hd__nor2_1
Xhold4380 _11809_/X vssd1 vssd1 vccd1 vccd1 _17093_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10145_ hold939/X hold3639/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__mux2_1
X_17810_ _17873_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4391 _17033_/Q vssd1 vssd1 vccd1 vccd1 hold4391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17741_ _17741_/CLK _17741_/D vssd1 vssd1 vccd1 vccd1 _17741_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3690 _17571_/Q vssd1 vssd1 vccd1 vccd1 hold3690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10076_ hold1801/X _16516_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__mux2_1
X_14953_ hold847/X _14952_/B _14952_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 hold848/A
+ sky130_fd_sc_hd__o211a_1
X_13904_ _15519_/A hold2276/X hold244/X vssd1 vssd1 vccd1 vccd1 _13905_/B sky130_fd_sc_hd__mux2_1
X_17672_ _17736_/CLK _17672_/D vssd1 vssd1 vccd1 vccd1 _17672_/Q sky130_fd_sc_hd__dfxtp_1
X_14884_ hold730/X _14894_/B vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__or2_1
X_16623_ _18192_/CLK _16623_/D vssd1 vssd1 vccd1 vccd1 _16623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _17732_/Q _13856_/B _13865_/C vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_23__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_23__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16554_ _18236_/CLK _16554_/D vssd1 vssd1 vccd1 vccd1 _16554_/Q sky130_fd_sc_hd__dfxtp_1
X_13766_ hold2111/X hold3273/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ hold3194/X _11171_/B _10977_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ _15521_/A hold1762/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15506_/B sky130_fd_sc_hd__mux2_1
X_12717_ _12777_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _17415_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16485_ _18398_/CLK _16485_/D vssd1 vssd1 vccd1 vccd1 _16485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13697_ hold1824/X hold3291/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13698_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18224_ _18224_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15436_ _17319_/Q _15479_/A2 _15446_/B1 hold259/X vssd1 vssd1 vccd1 vccd1 _15436_/X
+ sky130_fd_sc_hd__a22o_1
X_12648_ _12876_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _17392_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _18233_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
X_15367_ hold713/X _09357_/A _15484_/B1 hold703/X _15366_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/B sky130_fd_sc_hd__a221o_1
X_12579_ _12987_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _17369_/D sky130_fd_sc_hd__and2_1
X_17106_ _17268_/CLK _17106_/D vssd1 vssd1 vccd1 vccd1 _17106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _15105_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__or2_1
X_18086_ _18118_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ hold592/X _15484_/A2 _15451_/A2 hold578/X vssd1 vssd1 vccd1 vccd1 _15298_/X
+ sky130_fd_sc_hd__a22o_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _18073_/CLK _17037_/D vssd1 vssd1 vccd1 vccd1 _17037_/Q sky130_fd_sc_hd__dfxtp_1
X_14249_ hold1175/X _14266_/B _14248_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 fanout816/X vssd1 vssd1 vccd1 vccd1 _15208_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 fanout841/X vssd1 vssd1 vccd1 vccd1 _14813_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08810_ hold35/X hold471/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__mux2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ hold5717/X _10016_/B _09789_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09790_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _18374_/Q vssd1 vssd1 vccd1 vccd1 hold1006/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1017 _14235_/X vssd1 vssd1 vccd1 vccd1 _17918_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ hold41/X hold331/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__mux2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 _08300_/X vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ _18003_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1039 input39/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08672_ _09021_/A hold204/X vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09224_ _15553_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ hold2332/X _09164_/B _09154_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _09155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08106_ hold892/X hold919/X hold196/X vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_296_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17211_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ _14986_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08037_ _14330_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08037_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_225_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17873_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold840 hold840/A vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold851 input54/X vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold884 hold884/A vssd1 vssd1 vccd1 vccd1 hold884/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 hold895/A vssd1 vssd1 vccd1 vccd1 hold895/X sky130_fd_sc_hd__dlygate4sd3_1
X_09988_ _13078_/A _10016_/B _09987_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _16486_/D
+ sky130_fd_sc_hd__o211a_1
Xhold2230 _17902_/Q vssd1 vssd1 vccd1 vccd1 hold2230/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _17826_/Q vssd1 vssd1 vccd1 vccd1 hold2241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2252 _18098_/Q vssd1 vssd1 vccd1 vccd1 hold2252/X sky130_fd_sc_hd__dlygate4sd3_1
X_08939_ hold407/X hold612/X _08997_/S vssd1 vssd1 vccd1 vccd1 hold613/A sky130_fd_sc_hd__mux2_1
Xhold2263 _18305_/Q vssd1 vssd1 vccd1 vccd1 hold2263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2274 _18185_/Q vssd1 vssd1 vccd1 vccd1 hold2274/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1540 _18381_/Q vssd1 vssd1 vccd1 vccd1 hold1540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 _17937_/Q vssd1 vssd1 vccd1 vccd1 hold2285/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1551 _13056_/C vssd1 vssd1 vccd1 vccd1 hold1551/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2296 _08024_/X vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ hold3507/X _12362_/B _11949_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _11950_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1562 _13957_/X vssd1 vssd1 vccd1 vccd1 _17785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1573 _16312_/Q vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1584 _18429_/Q vssd1 vssd1 vccd1 vccd1 hold1584/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1595 _18277_/Q vssd1 vssd1 vccd1 vccd1 hold1595/X sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ hold2709/X hold3938/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ hold5106/X _13871_/B _11880_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _13710_/A _13620_/B vssd1 vssd1 vccd1 vccd1 _13620_/X sky130_fd_sc_hd__or2_1
X_10832_ hold1086/X hold5510/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _13776_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10763_ _17948_/Q _16745_/Q _10763_/S vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12502_ _17344_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16270_ _18431_/CLK _16270_/D vssd1 vssd1 vccd1 vccd1 _16270_/Q sky130_fd_sc_hd__dfxtp_1
X_13482_ _13674_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13482_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10694_ hold1175/X hold5254/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ _15221_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12433_ hold65/X hold520/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ hold2672/X hold609/X _15151_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _13873_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _12364_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ hold5965/X _14094_/B _14102_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 hold880/A
+ sky130_fd_sc_hd__o211a_1
X_11315_ hold1919/X hold3952/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__mux2_1
X_15083_ _15191_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12295_ _13822_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__nor2_1
X_14034_ _15541_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_5_7__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_11246_ hold1762/X hold3719/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11177_ _16883_/Q _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__and3_1
X_10128_ _10542_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10128_/X sky130_fd_sc_hd__or2_1
X_15985_ _17531_/CLK _15985_/D vssd1 vssd1 vccd1 vccd1 hold389/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17724_ _17724_/CLK _17724_/D vssd1 vssd1 vccd1 vccd1 _17724_/Q sky130_fd_sc_hd__dfxtp_1
X_10059_ _13270_/A _10380_/A _10058_/X vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__a21oi_1
X_14936_ _15205_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14936_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17877_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17655_ _17694_/CLK _17655_/D vssd1 vssd1 vccd1 vccd1 _17655_/Q sky130_fd_sc_hd__dfxtp_1
X_14867_ hold1555/X _14882_/B _14866_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14867_/X
+ sky130_fd_sc_hd__o211a_1
X_13818_ hold3764/X _13734_/A _13817_/X vssd1 vssd1 vccd1 vccd1 _13818_/Y sky130_fd_sc_hd__a21oi_1
X_16606_ _18222_/CLK _16606_/D vssd1 vssd1 vccd1 vccd1 _16606_/Q sky130_fd_sc_hd__dfxtp_1
X_17586_ _17749_/CLK _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ _15191_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _18095_/CLK _16537_/D vssd1 vssd1 vccd1 vccd1 _16537_/Q sky130_fd_sc_hd__dfxtp_1
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13749_/X sky130_fd_sc_hd__or2_1
XFILLER_0_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ _18381_/CLK _16468_/D vssd1 vssd1 vccd1 vccd1 _16468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15419_ hold550/X _15484_/A2 _15417_/X vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__a21o_1
X_18207_ _18267_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16399_ _18381_/CLK _16399_/D vssd1 vssd1 vccd1 vccd1 _16399_/Q sky130_fd_sc_hd__dfxtp_1
X_18138_ _18228_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5806 hold5934/X vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__buf_1
Xhold5817 hold5935/X vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5828 hold5828/A vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_12
Xhold114 hold264/X vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__clkbuf_8
Xhold5839 hold5839/A vssd1 vssd1 vccd1 vccd1 hold5839/X sky130_fd_sc_hd__clkbuf_4
Xhold125 hold317/X vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ _18069_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
Xhold136 hold2/X vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__buf_4
Xhold147 hold55/X vssd1 vssd1 vccd1 vccd1 input20/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold158 input34/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09911_ hold1006/X _16461_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__mux2_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 _09366_/Y vssd1 vssd1 vccd1 vccd1 _15484_/B1 sky130_fd_sc_hd__buf_6
Xfanout616 _09356_/Y vssd1 vssd1 vccd1 vccd1 _15446_/B1 sky130_fd_sc_hd__buf_6
Xfanout627 _09339_/Y vssd1 vssd1 vccd1 vccd1 _15481_/A1 sky130_fd_sc_hd__buf_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ hold2965/X hold4323/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__mux2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout638 _12849_/A vssd1 vssd1 vccd1 vccd1 _12825_/A sky130_fd_sc_hd__buf_4
Xfanout649 fanout660/X vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__buf_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ hold1610/X _16415_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__mux2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _09011_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _15983_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ hold359/X hold649/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__mux2_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ hold44/X hold310/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08587_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ hold1710/X _09218_/B _09206_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _09207_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _15521_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09069_ hold1075/X _09119_/A2 _09068_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _11658_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__or2_1
X_12080_ hold1231/X hold3347/X _12368_/C vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__mux2_1
Xhold670 hold670/A vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 hold681/A vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__buf_1
Xhold692 hold692/A vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11031_ _11031_/A _11031_/B vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__or2_1
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 _17878_/Q vssd1 vssd1 vccd1 vccd1 hold2060/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _14715_/X vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 _15760_/Q vssd1 vssd1 vccd1 vccd1 hold2082/X sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _17721_/CLK _15770_/D vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2093 _15814_/Q vssd1 vssd1 vccd1 vccd1 hold2093/X sky130_fd_sc_hd__dlygate4sd3_1
X_12982_ hold762/X _17505_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__mux2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 _15572_/Q vssd1 vssd1 vccd1 vccd1 hold1370/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1381 _16197_/Q vssd1 vssd1 vccd1 vccd1 hold1381/X sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ hold2268/X _14720_/B _14720_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14721_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ hold2040/X _17135_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__mux2_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _15160_/X vssd1 vssd1 vccd1 vccd1 _18363_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17456_/CLK _17440_/D vssd1 vssd1 vccd1 vccd1 _17440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _15099_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14652_/X sky130_fd_sc_hd__or2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ hold1603/X _17112_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__mux2_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ hold3291/X _13862_/B _13602_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _13603_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10815_ _11694_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__or2_1
X_17371_ _17981_/CLK _17371_/D vssd1 vssd1 vccd1 vccd1 _17371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ hold1438/X _14610_/B _14582_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14583_/X
+ sky130_fd_sc_hd__o211a_1
X_11795_ _17089_/Q _12341_/B _12341_/C vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16322_ _18460_/CLK _16322_/D vssd1 vssd1 vccd1 vccd1 _16322_/Q sky130_fd_sc_hd__dfxtp_1
X_13534_ hold4067/X _13829_/B _13533_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10746_ _11031_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_147_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18185_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16253_ _17447_/CLK _16253_/D vssd1 vssd1 vccd1 vccd1 _16253_/Q sky130_fd_sc_hd__dfxtp_1
X_13465_ hold5066/X _13859_/B _13464_/X _13753_/C1 vssd1 vssd1 vccd1 vccd1 _13465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _11136_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__or2_1
X_15204_ hold839/X _15221_/B _15203_/X _15070_/A vssd1 vssd1 vccd1 vccd1 hold840/A
+ sky130_fd_sc_hd__o211a_1
X_12416_ _12428_/A _12416_/B vssd1 vssd1 vccd1 vccd1 _17301_/D sky130_fd_sc_hd__and2_1
XFILLER_0_140_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16184_ _17482_/CLK _16184_/D vssd1 vssd1 vccd1 vccd1 _16184_/Q sky130_fd_sc_hd__dfxtp_1
X_13396_ hold4313/X _13886_/B _13395_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _13396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15135_ _15189_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__or2_1
X_12347_ _17273_/Q _12347_/B _13388_/S vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15066_ _15066_/A _15066_/B vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__and2_1
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ hold1422/X _17250_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__mux2_1
X_14017_ hold1201/X _14040_/B _14016_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14017_/X
+ sky130_fd_sc_hd__o211a_1
X_11229_ _12093_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15968_ _17323_/CLK _15968_/D vssd1 vssd1 vccd1 vccd1 hold559/A sky130_fd_sc_hd__dfxtp_1
X_17707_ _17734_/CLK _17707_/D vssd1 vssd1 vccd1 vccd1 _17707_/Q sky130_fd_sc_hd__dfxtp_1
X_14919_ hold2497/X _14946_/B _14918_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _14919_/X
+ sky130_fd_sc_hd__o211a_1
X_15899_ _17531_/CLK _15899_/D vssd1 vssd1 vccd1 vccd1 hold558/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08440_ hold2281/X _08440_/A2 _08439_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08440_/X
+ sky130_fd_sc_hd__o211a_1
X_17638_ _17734_/CLK _17638_/D vssd1 vssd1 vccd1 vccd1 _17638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ _08371_/A hold914/X vssd1 vssd1 vccd1 vccd1 _15817_/D sky130_fd_sc_hd__and2_1
X_17569_ _17731_/CLK _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5603 _09514_/X vssd1 vssd1 vccd1 vccd1 _16328_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5614 hold6026/X vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__buf_1
XFILLER_0_170_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5625 _16426_/Q vssd1 vssd1 vccd1 vccd1 hold5625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5636 _09634_/X vssd1 vssd1 vccd1 vccd1 _16368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4902 _10375_/X vssd1 vssd1 vccd1 vccd1 _16615_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5647 _16394_/Q vssd1 vssd1 vccd1 vccd1 hold5647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4913 _16514_/Q vssd1 vssd1 vccd1 vccd1 hold4913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5658 _10810_/X vssd1 vssd1 vccd1 vccd1 _16760_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4924 _12247_/X vssd1 vssd1 vccd1 vccd1 _17239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5669 _10927_/X vssd1 vssd1 vccd1 vccd1 _16799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4935 _17230_/Q vssd1 vssd1 vccd1 vccd1 hold4935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4946 _11992_/X vssd1 vssd1 vccd1 vccd1 _17154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4957 _16017_/Q vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4968 _11611_/X vssd1 vssd1 vccd1 vccd1 _17027_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout402 hold209/X vssd1 vssd1 vccd1 vccd1 _14433_/B sky130_fd_sc_hd__buf_6
Xhold4979 _16679_/Q vssd1 vssd1 vccd1 vccd1 hold4979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout413 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__buf_6
Xfanout424 _13998_/B vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__clkbuf_8
Xfanout435 _13808_/C vssd1 vssd1 vccd1 vccd1 _13805_/C sky130_fd_sc_hd__clkbuf_8
Xfanout446 fanout484/X vssd1 vssd1 vccd1 vccd1 _12353_/C sky130_fd_sc_hd__clkbuf_4
Xfanout457 fanout484/X vssd1 vssd1 vccd1 vccd1 _11171_/C sky130_fd_sc_hd__buf_4
X_09825_ _10779_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__or2_1
Xfanout468 _12368_/C vssd1 vssd1 vccd1 vccd1 _13844_/C sky130_fd_sc_hd__clkbuf_8
Xfanout479 _11672_/S vssd1 vssd1 vccd1 vccd1 _11792_/C sky130_fd_sc_hd__clkbuf_4
X_09756_ _09924_/A _09756_/B vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ hold8/X hold577/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__mux2_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09975_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__or2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _12438_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _15941_/D sky130_fd_sc_hd__and2_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _15491_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _15908_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ _11194_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10600_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _12051_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ hold4095/X _10643_/B _10530_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_240_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17649_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _17582_/Q _17116_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ hold5142/X _10558_/A2 _10461_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _13716_/A _12201_/B vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13181_ _13180_/X hold3179/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__mux2_1
X_10393_ hold4196/X _10589_/B _10392_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12132_ _12267_/A _12132_/B vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ _12255_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or2_1
X_16940_ _17852_/CLK _16940_/D vssd1 vssd1 vccd1 vccd1 _16940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11014_ hold3995/X _11210_/B _11013_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11014_/X
+ sky130_fd_sc_hd__o211a_1
X_16871_ _17981_/CLK _16871_/D vssd1 vssd1 vccd1 vccd1 _16871_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _17701_/CLK _15822_/D vssd1 vssd1 vccd1 vccd1 _15822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _17736_/CLK _15753_/D vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ hold3073/X _12964_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__mux2_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _12204_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__or2_1
X_14704_ _15205_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__or2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _17208_/CLK _15684_/D vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ hold3282/X _12895_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__mux2_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ hold2973/X _14666_/B _14634_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _14635_/X
+ sky130_fd_sc_hd__o211a_1
X_17423_ _17629_/CLK _17423_/D vssd1 vssd1 vccd1 vccd1 _17423_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _12243_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__or2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17516_/CLK _17354_/D vssd1 vssd1 vccd1 vccd1 _17354_/Q sky130_fd_sc_hd__dfxtp_1
X_14566_ _15492_/A _14573_/B hold934/X vssd1 vssd1 vccd1 vccd1 hold935/A sky130_fd_sc_hd__a21o_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ hold3781/X _12036_/A _11777_/X vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13517_ hold2182/X _17626_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__mux2_1
X_16305_ _17511_/CLK _16305_/D vssd1 vssd1 vccd1 vccd1 _16305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17285_ _17289_/CLK _17285_/D vssd1 vssd1 vccd1 vccd1 hold473/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ hold4625/X _11222_/B _10728_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14497_ _15231_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14497_/X sky130_fd_sc_hd__or2_1
X_16236_ _17754_/CLK _16236_/D vssd1 vssd1 vccd1 vccd1 _16236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13448_ _15840_/Q hold4220/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _17506_/CLK _16167_/D vssd1 vssd1 vccd1 vccd1 _16167_/Q sky130_fd_sc_hd__dfxtp_1
X_13379_ hold1445/X hold4200/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__mux2_1
Xhold4209 _16703_/Q vssd1 vssd1 vccd1 vccd1 hold4209/X sky130_fd_sc_hd__dlygate4sd3_1
X_15118_ hold5976/X _15113_/B hold430/X _15052_/A vssd1 vssd1 vccd1 vccd1 hold431/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16098_ _18414_/CLK _16098_/D vssd1 vssd1 vccd1 vccd1 _16098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3508 _11950_/X vssd1 vssd1 vccd1 vccd1 _17140_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3519 _17414_/Q vssd1 vssd1 vccd1 vccd1 hold3519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15049_ _15103_/A hold1970/X hold302/X vssd1 vssd1 vccd1 vccd1 _15050_/B sky130_fd_sc_hd__mux2_1
X_07940_ hold944/X _07988_/B vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__or2_1
Xhold2807 _18167_/Q vssd1 vssd1 vccd1 vccd1 hold2807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2818 _18372_/Q vssd1 vssd1 vccd1 vccd1 hold2818/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 _14516_/X vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07871_ _15549_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07871_/X sky130_fd_sc_hd__or2_1
X_09610_ hold5701/X _09992_/B _09609_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09610_/X
+ sky130_fd_sc_hd__o211a_1
X_09541_ hold5425/X _10025_/B _09540_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09541_/X
+ sky130_fd_sc_hd__o211a_1
X_09472_ _09472_/A _09472_/B _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09477_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_176_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ hold735/X _08445_/B vssd1 vssd1 vccd1 vccd1 _08423_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ hold949/X hold1087/X hold122/X vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ hold944/X _08335_/B vssd1 vssd1 vccd1 vccd1 _08285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5400 _09814_/X vssd1 vssd1 vccd1 vccd1 _16428_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5411 _16837_/Q vssd1 vssd1 vccd1 vccd1 hold5411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5422 _10888_/X vssd1 vssd1 vccd1 vccd1 _16786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5433 _16431_/Q vssd1 vssd1 vccd1 vccd1 hold5433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5444 _11293_/X vssd1 vssd1 vccd1 vccd1 _16921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5455 _09622_/X vssd1 vssd1 vccd1 vccd1 _16364_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4710 _17185_/Q vssd1 vssd1 vccd1 vccd1 hold4710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4721 _16852_/Q vssd1 vssd1 vccd1 vccd1 hold4721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5466 _17022_/Q vssd1 vssd1 vccd1 vccd1 hold5466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5477 _09697_/X vssd1 vssd1 vccd1 vccd1 _16389_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4732 _13681_/X vssd1 vssd1 vccd1 vccd1 _17680_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4743 _16685_/Q vssd1 vssd1 vccd1 vccd1 hold4743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5488 _16754_/Q vssd1 vssd1 vccd1 vccd1 hold5488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5499 _09547_/X vssd1 vssd1 vccd1 vccd1 _16339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4754 _09880_/X vssd1 vssd1 vccd1 vccd1 _16450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4765 _17141_/Q vssd1 vssd1 vccd1 vccd1 hold4765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4776 _13612_/X vssd1 vssd1 vccd1 vccd1 _17657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout210 _11150_/B vssd1 vssd1 vccd1 vccd1 _11156_/B sky130_fd_sc_hd__buf_4
Xfanout221 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10001_/B sky130_fd_sc_hd__buf_4
Xhold4787 _17659_/Q vssd1 vssd1 vccd1 vccd1 hold4787/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout232 _10610_/B vssd1 vssd1 vccd1 vccd1 _10580_/B sky130_fd_sc_hd__buf_2
Xhold4798 _11998_/X vssd1 vssd1 vccd1 vccd1 _17156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout243 _10649_/B vssd1 vssd1 vccd1 vccd1 _10640_/B sky130_fd_sc_hd__buf_4
Xfanout254 fanout299/X vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__clkbuf_4
Xfanout265 _11616_/A vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__buf_4
Xfanout276 fanout298/X vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__clkbuf_4
Xfanout287 _11688_/A vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__buf_4
X_09808_ hold5542/X _09998_/B _09807_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09808_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout298 fanout299/X vssd1 vssd1 vccd1 vccd1 fanout298/X sky130_fd_sc_hd__buf_4
X_09739_ hold4014/X _10025_/B _09738_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09739_/X
+ sky130_fd_sc_hd__o211a_1
X_12750_ _12753_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _17426_/D sky130_fd_sc_hd__and2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ hold4477/X _11798_/B _11700_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11701_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12876_/A _12681_/B vssd1 vssd1 vccd1 vccd1 _17403_/D sky130_fd_sc_hd__and2_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ hold2822/X _14433_/B _14419_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _14420_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ hold4303/X _11726_/B _11631_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14351_ hold826/X _17975_/Q hold275/X vssd1 vssd1 vccd1 vccd1 hold827/A sky130_fd_sc_hd__mux2_1
XFILLER_0_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ hold5342/X _11753_/B _11562_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13302_ _13302_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10514_ hold1326/X hold3338/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17070_ _17923_/CLK _17070_/D vssd1 vssd1 vccd1 vccd1 _17070_/Q sky130_fd_sc_hd__dfxtp_1
X_14282_ _15231_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11494_ hold3440/X _12323_/B _11493_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11494_/X
+ sky130_fd_sc_hd__o211a_1
X_16021_ _17523_/CLK _16021_/D vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__dfxtp_1
X_13233_ _13233_/A fanout2/A vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__and2_1
XFILLER_0_123_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ hold2183/X _16639_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ hold3129/X _13163_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__mux2_2
X_10376_ hold1469/X _16616_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ hold3366/X _12302_/B _12114_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12115_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17972_ _18069_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
X_13095_ _13183_/A1 _13093_/X _13094_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13095_/X
+ sky130_fd_sc_hd__o211a_1
X_12046_ hold3470/X _12347_/B _12045_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__o211a_1
X_16923_ _17908_/CLK _16923_/D vssd1 vssd1 vccd1 vccd1 _16923_/Q sky130_fd_sc_hd__dfxtp_1
X_16854_ _18059_/CLK _16854_/D vssd1 vssd1 vccd1 vccd1 _16854_/Q sky130_fd_sc_hd__dfxtp_1
X_15805_ _17748_/CLK _15805_/D vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13997_ hold1122/X _13986_/B _13996_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _13997_/X
+ sky130_fd_sc_hd__o211a_1
X_16785_ _18020_/CLK _16785_/D vssd1 vssd1 vccd1 vccd1 _16785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _17701_/CLK _15736_/D vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfxtp_1
X_12948_ _12951_/A _12948_/B vssd1 vssd1 vccd1 vccd1 _17492_/D sky130_fd_sc_hd__and2_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_162_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18455_ _18456_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
X_15667_ _17221_/CLK _15667_/D vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfxtp_1
X_12879_ _12885_/A _12879_/B vssd1 vssd1 vccd1 vccd1 _17469_/D sky130_fd_sc_hd__and2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17406_ _18458_/CLK _17406_/D vssd1 vssd1 vccd1 vccd1 _17406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14618_ _14726_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__or2_1
X_18386_ _18386_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _17266_/CLK _15598_/D vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17337_ _18417_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _17337_/Q sky130_fd_sc_hd__dfxtp_1
X_14549_ hold799/X _14553_/B vssd1 vssd1 vccd1 vccd1 _14549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08070_ _15529_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08070_/X sky130_fd_sc_hd__or2_1
X_17268_ _17268_/CLK _17268_/D vssd1 vssd1 vccd1 vccd1 _17268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16219_ _17453_/CLK _16219_/D vssd1 vssd1 vccd1 vccd1 _16219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17199_ _17263_/CLK _17199_/D vssd1 vssd1 vccd1 vccd1 _17199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4006 _16010_/Q vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4017 _10357_/X vssd1 vssd1 vccd1 vccd1 _16609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4028 _16347_/Q vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__buf_1
Xhold4039 _16839_/Q vssd1 vssd1 vccd1 vccd1 hold4039/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3305 _16666_/Q vssd1 vssd1 vccd1 vccd1 hold3305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3316 _11890_/X vssd1 vssd1 vccd1 vccd1 _17120_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08972_ _15491_/A _08972_/B vssd1 vssd1 vccd1 vccd1 _16103_/D sky130_fd_sc_hd__and2_1
Xhold3327 _10246_/X vssd1 vssd1 vccd1 vccd1 _16572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3338 _16662_/Q vssd1 vssd1 vccd1 vccd1 hold3338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3349 _16572_/Q vssd1 vssd1 vccd1 vccd1 hold3349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2604 _14837_/X vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 _14450_/X vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2626 _15648_/Q vssd1 vssd1 vccd1 vccd1 hold2626/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ hold1832/X _07924_/B _07922_/Y _08159_/A vssd1 vssd1 vccd1 vccd1 _07923_/X
+ sky130_fd_sc_hd__o211a_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__buf_4
Xhold2637 _15759_/Q vssd1 vssd1 vccd1 vccd1 hold2637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _15736_/Q vssd1 vssd1 vccd1 vccd1 hold2648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 _15659_/Q vssd1 vssd1 vccd1 vccd1 hold1903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _14015_/X vssd1 vssd1 vccd1 vccd1 _17813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 _16286_/Q vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1925 _18013_/Q vssd1 vssd1 vccd1 vccd1 hold1925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07854_ hold1370/X _07869_/B _07853_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07854_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1936 _17966_/Q vssd1 vssd1 vccd1 vccd1 hold1936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1947 _17780_/Q vssd1 vssd1 vccd1 vccd1 hold1947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1958 _15682_/Q vssd1 vssd1 vccd1 vccd1 hold1958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 _08097_/X vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07785_ _09438_/B vssd1 vssd1 vccd1 vccd1 _07785_/Y sky130_fd_sc_hd__inv_2
X_09524_ hold1379/X _13126_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__mux2_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09456_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09457_/C sky130_fd_sc_hd__or2_1
XFILLER_0_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ hold2513/X _08440_/A2 _08405_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _08406_/X
+ sky130_fd_sc_hd__o211a_1
X_09386_ _09386_/A _09386_/B _09392_/C _09386_/D vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08337_ hold624/X hold279/X vssd1 vssd1 vccd1 vccd1 _09399_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08268_ _15547_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08199_ _15533_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5230 _16333_/Q vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10230_ _10422_/A _10230_/B vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__or2_1
Xhold5241 _12331_/Y vssd1 vssd1 vccd1 vccd1 _17267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5252 _11184_/Y vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5263 _16729_/Q vssd1 vssd1 vccd1 vccd1 hold5263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5274 _11788_/Y vssd1 vssd1 vccd1 vccd1 _17086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4540 _16939_/Q vssd1 vssd1 vccd1 vccd1 hold4540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5285 _09996_/Y vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10161_ _10554_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10161_/X sky130_fd_sc_hd__or2_1
Xhold4551 _17256_/Q vssd1 vssd1 vccd1 vccd1 hold4551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5296 _11155_/Y vssd1 vssd1 vccd1 vccd1 _16875_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4562 _10333_/X vssd1 vssd1 vccd1 vccd1 _16601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4573 _16508_/Q vssd1 vssd1 vccd1 vccd1 hold4573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4584 _11704_/X vssd1 vssd1 vccd1 vccd1 _17058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4595 _17643_/Q vssd1 vssd1 vccd1 vccd1 hold4595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3850 _11181_/Y vssd1 vssd1 vccd1 vccd1 _11182_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3861 _16398_/Q vssd1 vssd1 vccd1 vccd1 hold3861/X sky130_fd_sc_hd__dlygate4sd3_1
X_10092_ _10380_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
Xhold3872 _11802_/Y vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3883 _17564_/Q vssd1 vssd1 vccd1 vccd1 hold3883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3894 _17572_/Q vssd1 vssd1 vccd1 vccd1 hold3894/X sky130_fd_sc_hd__dlygate4sd3_1
X_13920_ _14529_/A hold1683/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__mux2_1
X_13851_ hold3919/X _13779_/A _13850_/X vssd1 vssd1 vccd1 vccd1 _13851_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_5_22__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_22__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_12802_ hold1393/X hold3493/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16570_ _18224_/CLK _16570_/D vssd1 vssd1 vccd1 vccd1 _16570_/Q sky130_fd_sc_hd__dfxtp_1
X_13782_ _13791_/A _13782_/B vssd1 vssd1 vccd1 vccd1 _13782_/X sky130_fd_sc_hd__or2_1
X_10994_ hold2903/X hold4077/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__mux2_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ hold2087/X hold3077/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12733_/X sky130_fd_sc_hd__mux2_1
X_15521_ _15521_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _15489_/A _15452_/B _15452_/C _15452_/D vssd1 vssd1 vccd1 vccd1 _15452_/X
+ sky130_fd_sc_hd__or4_1
X_18240_ _18415_/CLK hold639/X vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ hold1985/X hold3022/X _12910_/S vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__mux2_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _15191_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ hold2042/X _17029_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15383_ _15481_/A1 _15375_/X _15382_/X _15481_/B1 hold5181/X vssd1 vssd1 vccd1 vccd1
+ _15383_/X sky130_fd_sc_hd__a32o_1
X_18171_ _18235_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12595_ hold2314/X hold3216/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17122_ _17282_/CLK _17122_/D vssd1 vssd1 vccd1 vccd1 _17122_/Q sky130_fd_sc_hd__dfxtp_1
X_14334_ _14728_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14334_/X sky130_fd_sc_hd__or2_1
X_11546_ hold1353/X _17006_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _17901_/CLK _17053_/D vssd1 vssd1 vccd1 vccd1 _17053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14265_ hold1463/X _14272_/B _14264_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11477_ hold1349/X hold5715/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__mux2_1
X_16004_ _18411_/CLK _16004_/D vssd1 vssd1 vccd1 vccd1 hold720/A sky130_fd_sc_hd__dfxtp_1
X_13216_ _13209_/X _13215_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17545_/D sky130_fd_sc_hd__o21a_1
X_10428_ _10524_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__or2_1
X_14196_ _15000_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13146_/X hold3156/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ _10551_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__or2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _18052_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
X_13078_ _13078_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__or2_1
X_12029_ hold1901/X _17167_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__mux2_1
X_16906_ _18432_/CLK _16906_/D vssd1 vssd1 vccd1 vccd1 _16906_/Q sky130_fd_sc_hd__dfxtp_1
X_17886_ _18051_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _18046_/CLK _16837_/D vssd1 vssd1 vccd1 vccd1 _16837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16768_ _18035_/CLK _16768_/D vssd1 vssd1 vccd1 vccd1 _16768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15719_ _17592_/CLK _15719_/D vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfxtp_1
X_16699_ _18225_/CLK _16699_/D vssd1 vssd1 vccd1 vccd1 _16699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ _12777_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _16231_/D sky130_fd_sc_hd__and2_1
X_18438_ _18438_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09171_ hold2348/X _09164_/B _09170_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09171_/X
+ sky130_fd_sc_hd__o211a_1
X_18369_ _18371_/CLK hold610/X vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ _15527_/A hold2630/X hold196/X vssd1 vssd1 vccd1 vccd1 _08123_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ hold906/X _08082_/B _08052_/X _08163_/A vssd1 vssd1 vccd1 vccd1 hold907/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3102 _17394_/Q vssd1 vssd1 vccd1 vccd1 hold3102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3113 _17448_/Q vssd1 vssd1 vccd1 vccd1 hold3113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3124 _17381_/Q vssd1 vssd1 vccd1 vccd1 hold3124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3135 _16534_/Q vssd1 vssd1 vccd1 vccd1 hold3135/X sky130_fd_sc_hd__buf_1
Xhold2401 _15851_/Q vssd1 vssd1 vccd1 vccd1 hold2401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3146 _10579_/Y vssd1 vssd1 vccd1 vccd1 _16683_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08955_ hold53/X _16095_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__mux2_1
Xhold2412 _08186_/X vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3157 _11742_/Y vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 _17106_/Q vssd1 vssd1 vccd1 vccd1 hold3168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 _17962_/Q vssd1 vssd1 vccd1 vccd1 hold2423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3179 _16531_/Q vssd1 vssd1 vccd1 vccd1 hold3179/X sky130_fd_sc_hd__buf_1
Xhold2434 _15019_/X vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2445 _18229_/Q vssd1 vssd1 vccd1 vccd1 hold2445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 _15867_/Q vssd1 vssd1 vccd1 vccd1 hold1700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 _09207_/X vssd1 vssd1 vccd1 vccd1 _16215_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07906_ _15529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__or2_1
Xhold2456 _17980_/Q vssd1 vssd1 vccd1 vccd1 hold2456/X sky130_fd_sc_hd__dlygate4sd3_1
X_08886_ hold126/X hold448/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__mux2_1
Xhold2467 _09306_/X vssd1 vssd1 vccd1 vccd1 _16263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1722 _17983_/Q vssd1 vssd1 vccd1 vccd1 hold1722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _18366_/Q vssd1 vssd1 vccd1 vccd1 hold2478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _14631_/X vssd1 vssd1 vccd1 vccd1 _18108_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1744 _17794_/Q vssd1 vssd1 vccd1 vccd1 hold1744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 _17970_/Q vssd1 vssd1 vccd1 vccd1 hold2489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1755 _14029_/X vssd1 vssd1 vccd1 vccd1 _17820_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1766 _08202_/X vssd1 vssd1 vccd1 vccd1 _15737_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07837_ _15515_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07837_/X sky130_fd_sc_hd__or2_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1777 _13031_/X vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _15880_/Q vssd1 vssd1 vccd1 vccd1 hold1788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1799 _17824_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09507_ _09903_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__or2_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09438_ _16305_/Q _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__or2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09369_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11400_ _12051_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12380_ _12380_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12425_/S sky130_fd_sc_hd__or2_2
XFILLER_0_118_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_70 hold784/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _15207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 _13252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _12018_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _15123_/A _14050_/B vssd1 vssd1 vccd1 vccd1 _14050_/X sky130_fd_sc_hd__or2_1
X_11262_ _12036_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_6__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5060 _17619_/Q vssd1 vssd1 vccd1 vccd1 hold5060/X sky130_fd_sc_hd__dlygate4sd3_1
X_13001_ hold3467/X _13000_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__mux2_1
X_10213_ hold4675/X _10619_/B _10212_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5071 _11428_/X vssd1 vssd1 vccd1 vccd1 _16966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5082 _17618_/Q vssd1 vssd1 vccd1 vccd1 hold5082/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5093 _13591_/X vssd1 vssd1 vccd1 vccd1 _17650_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11193_ hold3708/X _11097_/A _11192_/X vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4370 _11257_/X vssd1 vssd1 vccd1 vccd1 _16909_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10144_ hold4222/X _10589_/B _10143_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10144_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4381 _16640_/Q vssd1 vssd1 vccd1 vccd1 hold4381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4392 _11533_/X vssd1 vssd1 vccd1 vccd1 _17001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3680 _10609_/Y vssd1 vssd1 vccd1 vccd1 _16693_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17740_ _17740_/CLK _17740_/D vssd1 vssd1 vccd1 vccd1 _17740_/Q sky130_fd_sc_hd__dfxtp_1
X_10075_ _10588_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__nor2_1
Xhold3691 _13833_/Y vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14952_ _15221_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nand2_1
X_13903_ _13929_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _17759_/D sky130_fd_sc_hd__and2_1
Xhold2990 _07798_/X vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17671_ _17738_/CLK _17671_/D vssd1 vssd1 vccd1 vccd1 _17671_/Q sky130_fd_sc_hd__dfxtp_1
X_14883_ hold764/X _14882_/B _14882_/Y _14883_/C1 vssd1 vssd1 vccd1 vccd1 hold765/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16622_ _18266_/CLK _16622_/D vssd1 vssd1 vccd1 vccd1 _16622_/Q sky130_fd_sc_hd__dfxtp_1
X_13834_ _13864_/A _13834_/B vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _18319_/CLK _16553_/D vssd1 vssd1 vccd1 vccd1 _16553_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ hold5215/X _13859_/B _13764_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13765_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10977_ _11076_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or2_1
X_15504_ _15504_/A hold860/X vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12716_ hold3497/X _12715_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16484_ _18398_/CLK _16484_/D vssd1 vssd1 vccd1 vccd1 _16484_/Q sky130_fd_sc_hd__dfxtp_1
X_13696_ hold3539/X _13880_/B _13695_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18223_ _18223_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15435_ _15435_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__or2_1
X_12647_ hold2224/X _12646_/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15366_ _17340_/Q _15486_/B1 _15485_/B1 hold676/X vssd1 vssd1 vccd1 vccd1 _15366_/X
+ sky130_fd_sc_hd__a22o_1
X_18154_ _18224_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ hold3076/X _12577_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17105_ _17900_/CLK _17105_/D vssd1 vssd1 vccd1 vccd1 _17105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11529_ _11616_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__or2_1
X_14317_ hold2740/X _14326_/B _14316_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14317_/X
+ sky130_fd_sc_hd__o211a_1
X_18085_ _18149_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
X_15297_ hold512/X _09357_/A _15484_/B1 hold662/X _15296_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/B sky130_fd_sc_hd__a221o_1
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ _17852_/CLK _17036_/D vssd1 vssd1 vccd1 vccd1 _17036_/Q sky130_fd_sc_hd__dfxtp_1
X_14248_ _14517_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14248_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ hold1116/X _14202_/B _14178_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14179_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _15144_/C1 vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__buf_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _15491_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _15990_/D sky130_fd_sc_hd__and2_1
Xhold1007 _15184_/X vssd1 vssd1 vccd1 vccd1 _18374_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _17916_/Q vssd1 vssd1 vccd1 vccd1 hold1018/X sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ _18190_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1029 hold1069/X vssd1 vssd1 vccd1 vccd1 hold1070/A sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ hold35/X _15957_/Q _08727_/S vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17869_ _17891_/CLK hold749/X vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ hold1511/X _09216_/B _09222_/X _12843_/A vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _15537_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08105_ _15498_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _15691_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09085_ hold2752/X _09119_/A2 _09084_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09085_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08036_ hold1903/X _08033_/B _08035_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _08036_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold830 hold830/A vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 hold841/A vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold885 hold885/A vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 hold896/A vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_265_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__or2_1
Xhold2220 _15570_/Q vssd1 vssd1 vccd1 vccd1 hold2220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2231 _14199_/X vssd1 vssd1 vccd1 vccd1 _17902_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _15344_/A _08938_/B vssd1 vssd1 vccd1 vccd1 _16086_/D sky130_fd_sc_hd__and2_1
Xhold2242 _14041_/X vssd1 vssd1 vccd1 vccd1 _17826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2253 _14609_/X vssd1 vssd1 vccd1 vccd1 _18098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2264 _15625_/Q vssd1 vssd1 vccd1 vccd1 hold2264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1530 _15516_/X vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2275 _14791_/X vssd1 vssd1 vccd1 vccd1 _18185_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1541 _15198_/X vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 _14273_/X vssd1 vssd1 vccd1 vccd1 _17937_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _13033_/Y vssd1 vssd1 vccd1 vccd1 _17521_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ _12380_/B _08999_/B vssd1 vssd1 vccd1 vccd1 _08910_/S sky130_fd_sc_hd__or2_2
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2297 _17979_/Q vssd1 vssd1 vccd1 vccd1 hold2297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1563 _18049_/Q vssd1 vssd1 vccd1 vccd1 hold1563/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1574 _09417_/X vssd1 vssd1 vccd1 vccd1 _16294_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1585 hold6032/X vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__buf_1
X_10900_ hold4077/X _11210_/B _10899_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10900_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1596 _14983_/X vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ _13392_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__or2_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ hold5407/X _10897_/A2 _10830_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ hold1856/X _17637_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13551_/B sky130_fd_sc_hd__mux2_1
X_10762_ hold4371/X _10852_/A2 _10761_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _10762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12501_ hold44/X _12509_/A2 _12505_/A3 _12500_/X _09063_/A vssd1 vssd1 vccd1 vccd1
+ hold45/A sky130_fd_sc_hd__o311a_1
XFILLER_0_176_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13481_ hold2401/X hold4498/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_192_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10693_ hold3987/X _11747_/B _10692_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15220_ hold2693/X _15219_/B _15219_/Y _15030_/A vssd1 vssd1 vccd1 vccd1 _15220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _15344_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _17309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _15205_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__or2_1
X_12363_ hold3731/X _13392_/A _12362_/X vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__a21oi_1
X_14102_ hold799/X _14106_/B vssd1 vssd1 vccd1 vccd1 _14102_/X sky130_fd_sc_hd__or2_1
X_11314_ hold4403/X _11792_/B _11313_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__o211a_1
X_15082_ hold2932/X _15109_/B _15081_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15082_/X
+ sky130_fd_sc_hd__o211a_1
X_12294_ hold3165/X _12210_/A _12293_/X vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__a21oi_1
X_14033_ hold1167/X _14040_/B _14032_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14033_/X
+ sky130_fd_sc_hd__o211a_1
X_11245_ hold4455/X _11726_/B _11244_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _11245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11176_ _12331_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__nor2_1
X_10127_ hold1797/X hold3678/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__mux2_1
X_15984_ _17531_/CLK _15984_/D vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
X_17723_ _17723_/CLK _17723_/D vssd1 vssd1 vccd1 vccd1 _17723_/Q sky130_fd_sc_hd__dfxtp_1
X_14935_ hold822/X _14946_/B _14934_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 hold823/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10058_ _16510_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10058_/X sky130_fd_sc_hd__and3_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17654_ _17686_/CLK _17654_/D vssd1 vssd1 vccd1 vccd1 _17654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ _14866_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _18219_/CLK _16605_/D vssd1 vssd1 vccd1 vccd1 _16605_/Q sky130_fd_sc_hd__dfxtp_1
X_13817_ _17726_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13817_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17585_ _17745_/CLK _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
X_14797_ hold1706/X _14822_/B _14796_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14797_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18417_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16536_ _18126_/CLK _16536_/D vssd1 vssd1 vccd1 vccd1 _16536_/Q sky130_fd_sc_hd__dfxtp_1
X_13748_ hold1414/X hold3566/X _13844_/C vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16467_ _18386_/CLK _16467_/D vssd1 vssd1 vccd1 vccd1 _16467_/Q sky130_fd_sc_hd__dfxtp_1
X_13679_ hold1177/X hold4673/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18206_ _18206_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
X_15418_ hold551/X _09367_/A _15486_/B1 _17345_/Q vssd1 vssd1 vccd1 vccd1 _15418_/X
+ sky130_fd_sc_hd__a22o_1
X_16398_ _18424_/CLK _16398_/D vssd1 vssd1 vccd1 vccd1 _16398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _18230_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
X_15349_ hold530/X _09365_/B _09392_/C hold595/X _15348_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/C sky130_fd_sc_hd__a221o_1
Xhold5807 output95/X vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_12
Xhold5818 output72/X vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_12
Xhold104 hold64/X vssd1 vssd1 vccd1 vccd1 input23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5829 _18413_/Q vssd1 vssd1 vccd1 vccd1 hold5829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold319/X vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__clkbuf_4
X_18068_ _18070_/CLK hold744/X vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold148 input20/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ hold5405/X _10013_/B _09909_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09910_/X
+ sky130_fd_sc_hd__o211a_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _17855_/CLK _17019_/D vssd1 vssd1 vccd1 vccd1 _17019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 _09364_/Y vssd1 vssd1 vccd1 vccd1 _15451_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ hold5371/X _10025_/B _09840_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09841_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout617 _09356_/Y vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__clkbuf_4
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 hold816/X vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__clkbuf_8
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _12849_/A vssd1 vssd1 vccd1 vccd1 _12843_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ hold4329/X _11201_/B _09771_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09772_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ hold380/X hold527/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08654_ _12420_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _15949_/D sky130_fd_sc_hd__and2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _15916_/D sky130_fd_sc_hd__and2_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09206_ _15535_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09137_ hold2462/X _09177_/A2 _09136_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09137_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _15183_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _15533_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__or2_1
Xhold660 hold660/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 hold671/A vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11030_ hold1199/X hold4301/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11031_/B sky130_fd_sc_hd__mux2_1
Xhold682 hold682/A vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 hold693/A vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2050 _17901_/Q vssd1 vssd1 vccd1 vccd1 hold2050/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2061 _14149_/X vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _15569_/Q vssd1 vssd1 vccd1 vccd1 hold2072/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2083 _08251_/X vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12981_ _12987_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _17503_/D sky130_fd_sc_hd__and2_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2094 _18015_/Q vssd1 vssd1 vccd1 vccd1 hold2094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _07917_/X vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1371 _07854_/X vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ _14774_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__nand2_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ hold3353/X _12356_/B _11931_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11932_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1382 _09169_/X vssd1 vssd1 vccd1 vccd1 _16197_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _16213_/Q vssd1 vssd1 vccd1 vccd1 hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ hold4795/X _12341_/B _11862_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11863_/X
+ sky130_fd_sc_hd__o211a_1
X_14651_ hold2880/X _14666_/B _14650_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14651_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13767_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__or2_1
X_10814_ hold1412/X hold5574/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__mux2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17981_/CLK _17370_/D vssd1 vssd1 vccd1 vccd1 _17370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _15191_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__or2_1
X_11794_ _12343_/A _11794_/B vssd1 vssd1 vccd1 vccd1 _11794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ _18460_/CLK _16321_/D vssd1 vssd1 vccd1 vccd1 hold634/A sky130_fd_sc_hd__dfxtp_1
X_13533_ _13734_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _13533_/X sky130_fd_sc_hd__or2_1
X_10745_ hold2915/X hold5300/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13464_ _13758_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__or2_1
X_16252_ _17432_/CLK _16252_/D vssd1 vssd1 vccd1 vccd1 _16252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ hold1517/X hold3636/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15203_ hold747/X _15233_/B vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__or2_1
X_12415_ hold184/X hold474/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__mux2_1
X_13395_ _13749_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__or2_1
X_16183_ _17482_/CLK _16183_/D vssd1 vssd1 vccd1 vccd1 _16183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ hold1315/X _15161_/B _15133_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _15134_/X
+ sky130_fd_sc_hd__o211a_1
X_12346_ _13873_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_187_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18205_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15065_ _15227_/A hold2117/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15066_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_116_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18391_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12277_ hold4937/X _12377_/B _12276_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12277_/X
+ sky130_fd_sc_hd__o211a_1
X_14016_ hold949/X _14052_/B vssd1 vssd1 vccd1 vccd1 _14016_/X sky130_fd_sc_hd__or2_1
X_11228_ hold1767/X hold4815/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _16877_/Q _11735_/B _11735_/C vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15967_ _17313_/CLK _15967_/D vssd1 vssd1 vccd1 vccd1 hold701/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17706_ _17738_/CLK _17706_/D vssd1 vssd1 vccd1 vccd1 _17706_/Q sky130_fd_sc_hd__dfxtp_1
X_14918_ _14972_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14918_/X sky130_fd_sc_hd__or2_1
X_15898_ _17523_/CLK _15898_/D vssd1 vssd1 vccd1 vccd1 hold373/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17637_ _17701_/CLK _17637_/D vssd1 vssd1 vccd1 vccd1 _17637_/Q sky130_fd_sc_hd__dfxtp_1
X_14849_ hold1324/X _14882_/B _14848_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _15539_/A hold913/X hold122/X vssd1 vssd1 vccd1 vccd1 hold914/A sky130_fd_sc_hd__mux2_1
XFILLER_0_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17568_ _17728_/CLK _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ _18080_/CLK _16519_/D vssd1 vssd1 vccd1 vccd1 _16519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17499_ _18013_/CLK _17499_/D vssd1 vssd1 vccd1 vccd1 _17499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5604 _16947_/Q vssd1 vssd1 vccd1 vccd1 hold5604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5615 _16466_/Q vssd1 vssd1 vccd1 vccd1 hold5615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5626 _09712_/X vssd1 vssd1 vccd1 vccd1 _16394_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5637 _17201_/Q vssd1 vssd1 vccd1 vccd1 hold5637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4903 _17266_/Q vssd1 vssd1 vccd1 vccd1 hold4903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5648 _09616_/X vssd1 vssd1 vccd1 vccd1 _16362_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4914 _09976_/X vssd1 vssd1 vccd1 vccd1 _16482_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5659 _16890_/Q vssd1 vssd1 vccd1 vccd1 hold5659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4925 _17092_/Q vssd1 vssd1 vccd1 vccd1 hold4925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4936 _12124_/X vssd1 vssd1 vccd1 vccd1 _17198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4947 _16967_/Q vssd1 vssd1 vccd1 vccd1 hold4947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4958 _15481_/X vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4969 _17707_/Q vssd1 vssd1 vccd1 vccd1 hold4969/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout403 hold208/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__clkbuf_1
Xfanout414 _14162_/Y vssd1 vssd1 vccd1 vccd1 _14202_/B sky130_fd_sc_hd__clkbuf_8
Xfanout425 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13980_/B sky130_fd_sc_hd__buf_8
Xfanout436 _13808_/C vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__buf_6
Xfanout447 _11717_/C vssd1 vssd1 vccd1 vccd1 _12299_/C sky130_fd_sc_hd__clkbuf_8
X_09824_ hold2135/X _16432_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__mux2_1
Xfanout458 _13847_/C vssd1 vssd1 vccd1 vccd1 _13865_/C sky130_fd_sc_hd__clkbuf_8
Xfanout469 _12368_/C vssd1 vssd1 vccd1 vccd1 _12377_/C sky130_fd_sc_hd__clkbuf_8
X_09755_ hold2576/X hold4279/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09756_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08706_ _12428_/A hold93/X vssd1 vssd1 vccd1 vccd1 _15974_/D sky130_fd_sc_hd__and2_1
X_09686_ hold2942/X _16386_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ hold17/X hold238/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__mux2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ hold219/X hold715/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__mux2_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08499_ hold1146/X _08486_/B _08498_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _10548_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _11097_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
X_12200_ hold1519/X _17224_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_280_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18052_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13180_ hold3648/X _13179_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__mux2_2
X_10392_ _10551_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__or2_1
X_12131_ hold2707/X _17201_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12062_ hold1206/X hold4895/X _13388_/S vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__mux2_1
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__buf_8
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11013_ _11658_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11013_/X sky130_fd_sc_hd__or2_1
X_16870_ _18009_/CLK _16870_/D vssd1 vssd1 vccd1 vccd1 _16870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _17669_/CLK hold175/X vssd1 vssd1 vccd1 vccd1 _15821_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _17738_/CLK _15752_/D vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12964_ hold1752/X hold3059/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__mux2_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 _08308_/X vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ hold2832/X _14720_/B _14702_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14703_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ hold1497/X hold4769/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__mux2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _17779_/CLK hold838/X vssd1 vssd1 vccd1 vccd1 hold837/A sky130_fd_sc_hd__dfxtp_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ hold2228/X hold3121/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__mux2_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17428_/CLK _17422_/D vssd1 vssd1 vccd1 vccd1 _17422_/Q sky130_fd_sc_hd__dfxtp_1
X_14634_ _15189_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14634_/X sky130_fd_sc_hd__or2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ hold1025/X hold3168/X _12332_/C vssd1 vssd1 vccd1 vccd1 _11847_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17516_/CLK _17353_/D vssd1 vssd1 vccd1 vccd1 _17353_/Q sky130_fd_sc_hd__dfxtp_1
X_11777_ _17083_/Q _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _11777_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14565_ _15189_/A _14557_/Y hold1805/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16304_ _18460_/CLK hold618/X vssd1 vssd1 vccd1 vccd1 _16304_/Q sky130_fd_sc_hd__dfxtp_1
X_13516_ hold4889/X _13805_/B _13515_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__o211a_1
X_10728_ _11031_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
X_17284_ _17284_/CLK _17284_/D vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__dfxtp_1
X_14496_ hold1124/X _14487_/B _14495_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14496_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16235_ _17419_/CLK _16235_/D vssd1 vssd1 vccd1 vccd1 _16235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13447_ hold3963/X _13829_/B _13446_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _11637_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13378_ hold3390/X _13859_/B _13377_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__o211a_1
X_16166_ _17503_/CLK _16166_/D vssd1 vssd1 vccd1 vccd1 _16166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15117_ hold573/A _15125_/B vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__or2_1
X_12329_ _17267_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__and3_1
X_16097_ _17525_/CLK _16097_/D vssd1 vssd1 vccd1 vccd1 hold725/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3509 _17270_/Q vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__dlygate4sd3_1
X_15048_ _15058_/A _15048_/B vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2808 _14753_/X vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2819 _15178_/X vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07870_ hold2109/X _07865_/B _07869_/Y _12274_/C1 vssd1 vssd1 vccd1 vccd1 _07870_/X
+ sky130_fd_sc_hd__o211a_1
X_16999_ _17879_/CLK _16999_/D vssd1 vssd1 vccd1 vccd1 _16999_/Q sky130_fd_sc_hd__dfxtp_1
X_09540_ _09924_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_84_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17287_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18441_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09471_ _09472_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__or2_1
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08422_ hold1716/X _08433_/B _08421_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08353_ _09272_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__and2_1
XFILLER_0_176_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ hold816/X hold207/X vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__or2_4
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5401 _16495_/Q vssd1 vssd1 vccd1 vccd1 hold5401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5412 _10945_/X vssd1 vssd1 vccd1 vccd1 _16805_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5423 _16741_/Q vssd1 vssd1 vccd1 vccd1 hold5423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5434 _09727_/X vssd1 vssd1 vccd1 vccd1 _16399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4700 _16999_/Q vssd1 vssd1 vccd1 vccd1 hold4700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5445 _16778_/Q vssd1 vssd1 vccd1 vccd1 hold5445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4711 _11989_/X vssd1 vssd1 vccd1 vccd1 _17153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5456 _16989_/Q vssd1 vssd1 vccd1 vccd1 hold5456/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5467 _11500_/X vssd1 vssd1 vccd1 vccd1 _16990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4722 _10990_/X vssd1 vssd1 vccd1 vccd1 _16820_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4733 _17248_/Q vssd1 vssd1 vccd1 vccd1 hold4733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5478 _16862_/Q vssd1 vssd1 vccd1 vccd1 hold5478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4744 _10489_/X vssd1 vssd1 vccd1 vccd1 _16653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5489 _10696_/X vssd1 vssd1 vccd1 vccd1 _16722_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4755 _17734_/Q vssd1 vssd1 vccd1 vccd1 hold4755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4766 _11857_/X vssd1 vssd1 vccd1 vccd1 _17109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout200 _11210_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__buf_4
Xhold4777 _16549_/Q vssd1 vssd1 vccd1 vccd1 hold4777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4788 _13522_/X vssd1 vssd1 vccd1 vccd1 _17627_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout211 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _11150_/B sky130_fd_sc_hd__buf_4
XFILLER_0_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout222 _10558_/A2 vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__buf_4
Xfanout233 _10465_/A2 vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__clkbuf_4
Xhold4799 _16624_/Q vssd1 vssd1 vccd1 vccd1 hold4799/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout244 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__buf_4
Xfanout255 _13674_/A vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout266 fanout299/X vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__buf_4
Xfanout277 _12243_/A vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__buf_4
X_09807_ _09903_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__or2_1
Xfanout288 fanout298/X vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__buf_2
X_07999_ _14740_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _07999_/X sky130_fd_sc_hd__or2_1
Xfanout299 _09493_/Y vssd1 vssd1 vccd1 vccd1 fanout299/X sky130_fd_sc_hd__clkbuf_8
Xclkbuf_5_21__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_21__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_09738_ _09924_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _09975_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__or2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _12153_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _17403_/Q hold2214/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__mux2_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__or2_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11562_ _11658_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__or2_1
X_14350_ _14350_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _17974_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ hold4387/X _10631_/B _10512_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10513_/X
+ sky130_fd_sc_hd__o211a_1
X_13301_ _13300_/X hold3699/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ hold2429/X _14266_/B _14280_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ _11649_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13232_ _13225_/X _13231_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__o21a_1
X_16020_ _17528_/CLK _16020_/D vssd1 vssd1 vccd1 vccd1 hold692/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ hold5582/X _10897_/A2 _10443_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13163_ _13162_/X hold3645/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ hold4901/X _10465_/A2 _10374_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _10375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ _12210_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17971_ _18003_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
X_13094_ _13094_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__or2_1
Xhold5990 _17348_/Q vssd1 vssd1 vccd1 vccd1 hold5990/X sky130_fd_sc_hd__dlygate4sd3_1
X_12045_ _12243_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__or2_1
X_16922_ _17898_/CLK _16922_/D vssd1 vssd1 vccd1 vccd1 _16922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ _18066_/CLK _16853_/D vssd1 vssd1 vccd1 vccd1 _16853_/Q sky130_fd_sc_hd__dfxtp_1
X_15804_ _17737_/CLK _15804_/D vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfxtp_1
X_16784_ _18052_/CLK _16784_/D vssd1 vssd1 vccd1 vccd1 _16784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _15123_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13996_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15735_ _17738_/CLK _15735_/D vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ hold3380/X _12946_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18454_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
X_15666_ _17592_/CLK hold907/X vssd1 vssd1 vccd1 vccd1 hold906/A sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ hold3258/X _12877_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _18456_/CLK _17405_/D vssd1 vssd1 vccd1 vccd1 _17405_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ hold1505/X _14610_/B _14616_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14617_/X
+ sky130_fd_sc_hd__o211a_1
X_11829_ _13797_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__or2_1
X_18385_ _18385_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_15597_ _17170_/CLK _15597_/D vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336_ _18417_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _17336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ hold1911/X _14541_/B _14547_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14548_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_131_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18381_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17267_ _17865_/CLK _17267_/D vssd1 vssd1 vccd1 vccd1 _17267_/Q sky130_fd_sc_hd__dfxtp_1
X_14479_ _15105_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16218_ _17453_/CLK _16218_/D vssd1 vssd1 vccd1 vccd1 _16218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17198_ _17275_/CLK _17198_/D vssd1 vssd1 vccd1 vccd1 _17198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4007 _15413_/X vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4018 _16630_/Q vssd1 vssd1 vccd1 vccd1 hold4018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _17494_/CLK _16149_/D vssd1 vssd1 vccd1 vccd1 _16149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4029 _10050_/Y vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3306 _10432_/X vssd1 vssd1 vccd1 vccd1 _16634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3317 _17361_/Q vssd1 vssd1 vccd1 vccd1 hold3317/X sky130_fd_sc_hd__dlygate4sd3_1
X_08971_ hold219/X hold717/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__mux2_1
Xhold3328 _16414_/Q vssd1 vssd1 vccd1 vccd1 hold3328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3339 _10420_/X vssd1 vssd1 vccd1 vccd1 _16630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2605 _16210_/Q vssd1 vssd1 vccd1 vccd1 hold2605/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _15545_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__nand2_1
Xhold2616 _17819_/Q vssd1 vssd1 vccd1 vccd1 hold2616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2627 _08014_/X vssd1 vssd1 vccd1 vccd1 _15648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 _08249_/X vssd1 vssd1 vccd1 vccd1 _15759_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 _08200_/X vssd1 vssd1 vccd1 vccd1 _15736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _08036_/X vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1915 _07803_/Y vssd1 vssd1 vccd1 vccd1 hold1915/X sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _14866_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__or2_1
Xhold1926 _14430_/X vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1937 _14333_/X vssd1 vssd1 vccd1 vccd1 _17966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1948 _15571_/Q vssd1 vssd1 vccd1 vccd1 hold1948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 _08085_/X vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _18461_/Q vssd1 vssd1 vccd1 vccd1 _14556_/A sky130_fd_sc_hd__inv_2
XFILLER_0_190_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09523_ hold3831/X _10001_/B _09522_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09523_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09454_ _09455_/B _09481_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _16311_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08405_ _15519_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09385_ hold5845/A _09342_/B _09342_/Y _09384_/X _12442_/A vssd1 vssd1 vccd1 vccd1
+ _09385_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_219_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17799_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08336_ hold1971/X _08336_/A2 _08335_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ hold1850/X _08268_/B _08266_/Y _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08198_ hold1282/X _08209_/B _08197_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08198_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5220 _15433_/X vssd1 vssd1 vccd1 vccd1 _15434_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_5_5__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
Xhold5231 _10008_/Y vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5242 _16337_/Q vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5253 _11185_/Y vssd1 vssd1 vccd1 vccd1 _16885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5264 _11196_/Y vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4530 _17279_/Q vssd1 vssd1 vccd1 vccd1 hold4530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5275 _16330_/Q vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10160_ hold1505/X hold3728/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__mux2_1
Xhold5286 _09997_/Y vssd1 vssd1 vccd1 vccd1 _16489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4541 _11251_/X vssd1 vssd1 vccd1 vccd1 _16907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4552 _12202_/X vssd1 vssd1 vccd1 vccd1 _17224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5297 _16730_/Q vssd1 vssd1 vccd1 vccd1 hold5297/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4563 _17662_/Q vssd1 vssd1 vccd1 vccd1 hold4563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4574 _09958_/X vssd1 vssd1 vccd1 vccd1 _16476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3840 _10063_/Y vssd1 vssd1 vccd1 vccd1 _16511_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4585 _16955_/Q vssd1 vssd1 vccd1 vccd1 hold4585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4596 _13474_/X vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3851 _11182_/Y vssd1 vssd1 vccd1 vccd1 _16884_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10091_ hold1783/X hold3662/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__mux2_1
Xhold3862 _09628_/X vssd1 vssd1 vccd1 vccd1 _16366_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3873 _11803_/Y vssd1 vssd1 vccd1 vccd1 _17091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3884 _13812_/Y vssd1 vssd1 vccd1 vccd1 _13813_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3895 _13836_/Y vssd1 vssd1 vccd1 vccd1 _13837_/B sky130_fd_sc_hd__dlygate4sd3_1
X_13850_ _17737_/Q _13880_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12801_ _12804_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _17443_/D sky130_fd_sc_hd__and2_1
X_13781_ hold2216/X _17714_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__mux2_1
X_10993_ hold5534/X _11216_/B _10992_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ hold2557/X _15560_/A2 _15519_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _15520_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12756_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _17420_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ hold151/X _15451_/A2 _15484_/B1 hold557/X _15446_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/D sky130_fd_sc_hd__a221o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _15502_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _17397_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ hold2887/X hold209/X _14401_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _14402_/X
+ sky130_fd_sc_hd__o211a_1
X_11614_ hold4627/X _12320_/B _11613_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11614_/X
+ sky130_fd_sc_hd__o211a_1
X_18170_ _18228_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_15382_ _15471_/A _15382_/B _15382_/C _15382_/D vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_93_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ _15506_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _17374_/D sky130_fd_sc_hd__and2_1
X_17121_ _17281_/CLK _17121_/D vssd1 vssd1 vccd1 vccd1 _17121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14333_ hold1936/X _14333_/A2 _14332_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14333_/X
+ sky130_fd_sc_hd__o211a_1
X_11545_ hold4289/X _11735_/B _11544_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _17902_/CLK _17052_/D vssd1 vssd1 vccd1 vccd1 _17052_/Q sky130_fd_sc_hd__dfxtp_1
X_11476_ hold5707/X _11762_/B _11475_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11476_/X
+ sky130_fd_sc_hd__o211a_1
X_14264_ _15105_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__or2_1
X_16003_ _18410_/CLK _16003_/D vssd1 vssd1 vccd1 vccd1 hold687/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13215_ _13311_/A1 _13213_/X _13214_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13215_/X
+ sky130_fd_sc_hd__o211a_1
X_10427_ hold1565/X hold4561/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14195_ hold5970/X _14198_/B hold467/X _13933_/A vssd1 vssd1 vccd1 vccd1 hold468/A
+ sky130_fd_sc_hd__o211a_1
X_10358_ hold2612/X _16610_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__mux2_1
X_13146_ _17569_/Q _17103_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _18020_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
X_13077_ _13076_/X hold3545/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__mux2_1
X_10289_ hold2868/X _16587_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__mux2_1
X_12028_ hold3400/X _12314_/B _12027_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12028_/X
+ sky130_fd_sc_hd__o211a_1
X_16905_ _18431_/CLK _16905_/D vssd1 vssd1 vccd1 vccd1 _16905_/Q sky130_fd_sc_hd__dfxtp_1
X_17885_ _18073_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16836_ _18305_/CLK _16836_/D vssd1 vssd1 vccd1 vccd1 _16836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _18190_/CLK _16767_/D vssd1 vssd1 vccd1 vccd1 _16767_/Q sky130_fd_sc_hd__dfxtp_1
X_13979_ hold1065/X _13986_/B _13978_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _13979_/X
+ sky130_fd_sc_hd__o211a_1
X_15718_ _17253_/CLK _15718_/D vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfxtp_1
X_16698_ _18192_/CLK _16698_/D vssd1 vssd1 vccd1 vccd1 _16698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _18438_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_312_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17724_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15649_ _17257_/CLK _15649_/D vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ _15553_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__or2_1
X_18368_ _18422_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ _13931_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__and2_1
X_17319_ _17345_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 _17319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _18315_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
X_08052_ hold892/X _08094_/B vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3103 _17397_/Q vssd1 vssd1 vccd1 vccd1 hold3103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3114 _12815_/X vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3125 _12614_/X vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3136 _10611_/Y vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2402 _08442_/X vssd1 vssd1 vccd1 vccd1 _15851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3147 _17120_/Q vssd1 vssd1 vccd1 vccd1 hold3147/X sky130_fd_sc_hd__dlygate4sd3_1
X_08954_ _15473_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _16094_/D sky130_fd_sc_hd__and2_1
Xhold3158 _11743_/Y vssd1 vssd1 vccd1 vccd1 _17071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2413 _17373_/Q vssd1 vssd1 vccd1 vccd1 hold2413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3169 _12327_/Y vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _14325_/X vssd1 vssd1 vccd1 vccd1 _17962_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 _15859_/Q vssd1 vssd1 vccd1 vccd1 hold2435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 _14881_/X vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07905_ hold2622/X _07918_/B _07904_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07905_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1701 _08477_/X vssd1 vssd1 vccd1 vccd1 _15867_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1712 _15600_/Q vssd1 vssd1 vccd1 vccd1 hold1712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 _16184_/Q vssd1 vssd1 vccd1 vccd1 hold2457/X sky130_fd_sc_hd__dlygate4sd3_1
X_08885_ _15314_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _16060_/D sky130_fd_sc_hd__and2_1
Xhold1723 _18111_/Q vssd1 vssd1 vccd1 vccd1 hold1723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 _15699_/Q vssd1 vssd1 vccd1 vccd1 hold2468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _17872_/Q vssd1 vssd1 vccd1 vccd1 hold1734/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2479 _15166_/X vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 _13975_/X vssd1 vssd1 vccd1 vccd1 _17794_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07836_ hold2256/X _07865_/B _07835_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07836_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1756 _16318_/Q vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1767 _18426_/Q vssd1 vssd1 vccd1 vccd1 hold1767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1778 _18009_/Q vssd1 vssd1 vccd1 vccd1 hold1778/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1789 _08506_/X vssd1 vssd1 vccd1 vccd1 _15880_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_154_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09506_ hold1927/X _16326_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _07804_/A _09483_/A _15314_/A hold617/X vssd1 vssd1 vccd1 vccd1 hold618/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _09386_/B _09369_/B _09369_/C _09369_/D vssd1 vssd1 vccd1 vccd1 _09368_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _15543_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ _15521_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_60 hold173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_71 hold799/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_82 _15207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11330_ hold1229/X _16934_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__mux2_1
XANTENNA_93 _14286_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ hold894/X hold3156/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11262_/B sky130_fd_sc_hd__mux2_1
Xhold5050 _16857_/Q vssd1 vssd1 vccd1 vccd1 hold5050/X sky130_fd_sc_hd__dlygate4sd3_1
X_10212_ _10524_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__or2_1
Xhold5061 _13402_/X vssd1 vssd1 vccd1 vccd1 _17587_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13000_ hold2288/X _07826_/A _13000_/S vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5072 _16474_/Q vssd1 vssd1 vccd1 vccd1 hold5072/X sky130_fd_sc_hd__dlygate4sd3_1
X_11192_ _16888_/Q _11192_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__and3_1
Xhold5083 _13399_/X vssd1 vssd1 vccd1 vccd1 _17586_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5094 _16551_/Q vssd1 vssd1 vccd1 vccd1 hold5094/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4360 _10162_/X vssd1 vssd1 vccd1 vccd1 _16544_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10143_ _10551_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__or2_1
Xhold4371 _16776_/Q vssd1 vssd1 vccd1 vccd1 hold4371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4382 _10354_/X vssd1 vssd1 vccd1 vccd1 _16608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4393 _17226_/Q vssd1 vssd1 vccd1 vccd1 hold4393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3670 _17730_/Q vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14951_ hold1103/X _14946_/B _14950_/Y _15070_/A vssd1 vssd1 vccd1 vccd1 _14951_/X
+ sky130_fd_sc_hd__o211a_1
X_10074_ _13310_/A _10506_/A _10073_/X vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__a21oi_1
Xhold3681 _16344_/Q vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3692 _13834_/Y vssd1 vssd1 vccd1 vccd1 _17731_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13902_ _14511_/A hold894/X hold244/X vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2980 _08455_/X vssd1 vssd1 vccd1 vccd1 _15856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17670_ _17734_/CLK _17670_/D vssd1 vssd1 vccd1 vccd1 _17670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _15221_/A _14882_/B vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__nand2_1
Xhold2991 _07799_/Y vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16621_ _18266_/CLK _16621_/D vssd1 vssd1 vccd1 vccd1 _16621_/Q sky130_fd_sc_hd__dfxtp_1
X_13833_ hold3690/X _13737_/A _13832_/X vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16552_ _18205_/CLK _16552_/D vssd1 vssd1 vccd1 vccd1 _16552_/Q sky130_fd_sc_hd__dfxtp_1
X_13764_ _13764_/A _13764_/B vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__or2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ hold2361/X _16816_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ hold826/X _18431_/Q _15505_/S vssd1 vssd1 vccd1 vccd1 hold860/A sky130_fd_sc_hd__mux2_1
X_12715_ hold2541/X hold3489/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16483_ _18388_/CLK _16483_/D vssd1 vssd1 vccd1 vccd1 _16483_/Q sky130_fd_sc_hd__dfxtp_1
X_13695_ _13791_/A _13695_/B vssd1 vssd1 vccd1 vccd1 _13695_/X sky130_fd_sc_hd__or2_1
X_18222_ _18222_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _15473_/A _15434_/B vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__and2_1
X_12646_ hold1346/X _17393_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _18268_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
X_15365_ hold469/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ hold2483/X hold3071/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _17908_/CLK _17104_/D vssd1 vssd1 vccd1 vccd1 _17104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _15103_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__or2_1
X_18084_ _18265_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ hold1322/X _17000_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__mux2_1
X_15296_ _17333_/Q _09362_/C _15485_/B1 hold472/X vssd1 vssd1 vccd1 vccd1 _15296_/X
+ sky130_fd_sc_hd__a22o_1
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 input35/X vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17035_ _17884_/CLK _17035_/D vssd1 vssd1 vccd1 vccd1 _17035_/Q sky130_fd_sc_hd__dfxtp_1
X_14247_ hold2809/X _14266_/B _14246_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14247_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11459_ hold2197/X hold4137/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14178_ _14517_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14178_/X sky130_fd_sc_hd__or2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13129_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__and2_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _15565_/Q vssd1 vssd1 vccd1 vccd1 hold1008/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _18025_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1019 _14229_/X vssd1 vssd1 vccd1 vccd1 _17916_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _12420_/A hold417/X vssd1 vssd1 vccd1 vccd1 _15956_/D sky130_fd_sc_hd__and2_1
X_17868_ _17900_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16819_ _18054_/CLK _16819_/D vssd1 vssd1 vccd1 vccd1 _16819_/Q sky130_fd_sc_hd__dfxtp_1
X_17799_ _17799_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _15551_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ hold1742/X _09164_/B _09152_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _09153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ _14218_/A hold2840/X hold196/X vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _14984_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08035_ _15549_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08035_/X sky130_fd_sc_hd__or2_1
Xhold820 hold820/A vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 hold831/A vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold864 hold864/A vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold886 hold886/A vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 becStatus[2] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ hold2518/X hold5512/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__mux2_1
Xhold2210 hold2210/A vssd1 vssd1 vccd1 vccd1 input69/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2221 _07850_/X vssd1 vssd1 vccd1 vccd1 _15570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 _18293_/Q vssd1 vssd1 vccd1 vccd1 hold2232/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ hold68/X hold396/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08938_/B sky130_fd_sc_hd__mux2_1
Xhold2243 _15714_/Q vssd1 vssd1 vccd1 vccd1 hold2243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2254 _15586_/Q vssd1 vssd1 vccd1 vccd1 hold2254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1520 _07929_/X vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2265 _07965_/X vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 _18218_/Q vssd1 vssd1 vccd1 vccd1 hold1531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 _17760_/Q vssd1 vssd1 vccd1 vccd1 hold2276/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2287 _17993_/Q vssd1 vssd1 vccd1 vccd1 hold2287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _17951_/Q vssd1 vssd1 vccd1 vccd1 hold1542/X sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ _17520_/Q _08868_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__or3b_4
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1553 _17959_/Q vssd1 vssd1 vccd1 vccd1 hold1553/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2298 _17964_/Q vssd1 vssd1 vccd1 vccd1 hold2298/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _14506_/X vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1575 _16241_/Q vssd1 vssd1 vccd1 vccd1 hold1575/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1586 _09409_/X vssd1 vssd1 vccd1 vccd1 _16290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_234_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17283_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07819_ _15559_/A _15231_/A vssd1 vssd1 vccd1 vccd1 _09495_/C sky130_fd_sc_hd__nand2_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _18088_/Q vssd1 vssd1 vccd1 vccd1 hold1597/X sky130_fd_sc_hd__dlygate4sd3_1
X_08799_ hold68/X hold707/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold708/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _11103_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _11631_/A _10761_/B vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12500_ _17343_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ hold4395/X _13832_/B _13479_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13480_/X
+ sky130_fd_sc_hd__o211a_1
X_10692_ _11652_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ hold50/X hold293/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ hold806/X _15161_/B _15149_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 hold807/A
+ sky130_fd_sc_hd__o211a_1
X_12362_ _17278_/Q _12362_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ hold2236/X _14105_/A2 _14100_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _11697_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15081_ _15189_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__or2_1
X_12293_ _17255_/Q _12302_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ _15105_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__or2_1
X_11244_ _11631_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ hold5254/X _11658_/A _11174_/X vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4190 _16556_/Q vssd1 vssd1 vccd1 vccd1 hold4190/X sky130_fd_sc_hd__dlygate4sd3_1
X_10126_ hold4165/X _10589_/B _10125_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _17345_/CLK _15983_/D vssd1 vssd1 vccd1 vccd1 hold527/A sky130_fd_sc_hd__dfxtp_1
X_17722_ _17722_/CLK _17722_/D vssd1 vssd1 vccd1 vccd1 _17722_/Q sky130_fd_sc_hd__dfxtp_1
X_10057_ _10588_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__nor2_1
X_14934_ hold747/X _14962_/B vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _17749_/CLK _17653_/D vssd1 vssd1 vccd1 vccd1 _17653_/Q sky130_fd_sc_hd__dfxtp_1
X_14865_ hold2283/X _14880_/B _14864_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14865_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_188_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16604_ _18226_/CLK _16604_/D vssd1 vssd1 vccd1 vccd1 _16604_/Q sky130_fd_sc_hd__dfxtp_1
X_13816_ _13822_/A _13816_/B vssd1 vssd1 vccd1 vccd1 _13816_/Y sky130_fd_sc_hd__nor2_1
X_17584_ _17584_/CLK _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14796_ _14850_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14796_/X sky130_fd_sc_hd__or2_1
X_16535_ _18221_/CLK _16535_/D vssd1 vssd1 vccd1 vccd1 _16535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ hold4755/X _13859_/B _13746_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13747_/X
+ sky130_fd_sc_hd__o211a_1
X_10959_ _11061_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__or2_1
X_16466_ _18373_/CLK _16466_/D vssd1 vssd1 vccd1 vccd1 _16466_/Q sky130_fd_sc_hd__dfxtp_1
X_13678_ hold4848/X _13856_/B _13677_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13678_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18205_ _18205_/CLK hold961/X vssd1 vssd1 vccd1 vccd1 hold960/A sky130_fd_sc_hd__dfxtp_1
X_15417_ hold495/X _09392_/B _09392_/C hold323/X vssd1 vssd1 vccd1 vccd1 _15417_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12629_ hold3086/X _12628_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__mux2_1
X_16397_ _18420_/CLK _16397_/D vssd1 vssd1 vccd1 vccd1 _16397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18136_ _18220_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18050_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ hold554/X _09386_/A _15451_/A2 hold561/X vssd1 vssd1 vccd1 vccd1 _15348_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5808 hold5932/X vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5819 _18403_/Q vssd1 vssd1 vccd1 vccd1 hold5819/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 input23/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__buf_1
X_18067_ _18067_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
X_15279_ hold239/X _15485_/A2 _15447_/B1 hold165/X _15278_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold56/X vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__buf_4
XFILLER_0_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17018_ _17898_/CLK _17018_/D vssd1 vssd1 vccd1 vccd1 _17018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09840_ _09924_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__or2_1
Xfanout607 _09364_/Y vssd1 vssd1 vccd1 vccd1 _09392_/D sky130_fd_sc_hd__buf_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout618 _09354_/Y vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__buf_6
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout629 hold815/X vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__buf_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _11082_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__or2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08722_ _12428_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _15982_/D sky130_fd_sc_hd__and2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08653_ hold44/X hold414/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ hold65/X hold569/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ hold2520/X _09218_/B _09204_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _09205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09136_ _15519_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__or2_1
X_09067_ _15182_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__or2_2
XFILLER_0_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08018_ hold1105/X _08029_/B _08017_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _08018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold650 hold650/A vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 hold661/A vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 hold672/A vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold683 hold683/A vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold694/A vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ _10491_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__or2_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2040 _15675_/Q vssd1 vssd1 vccd1 vccd1 hold2040/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 _14197_/X vssd1 vssd1 vccd1 vccd1 _17901_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2062 _18451_/Q vssd1 vssd1 vccd1 vccd1 hold2062/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2073 _07848_/X vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12980_ hold3100/X _12979_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__mux2_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2084 _15705_/Q vssd1 vssd1 vccd1 vccd1 hold2084/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 _14051_/X vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2095 _14434_/X vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _16209_/Q vssd1 vssd1 vccd1 vccd1 hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 _16231_/Q vssd1 vssd1 vccd1 vccd1 hold1372/X sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ _12267_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__or2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 _17818_/Q vssd1 vssd1 vccd1 vccd1 hold1383/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _09203_/X vssd1 vssd1 vccd1 vccd1 _16213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _15205_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__or2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _12246_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11862_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ hold1189/X _17654_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__mux2_1
X_10813_ hold4716/X _11192_/B _10812_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ hold2893/X _14612_/B _14580_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14581_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ hold3713/X _11697_/A _11792_/X vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _18460_/CLK _16320_/D vssd1 vssd1 vccd1 vccd1 _16320_/Q sky130_fd_sc_hd__dfxtp_1
X_13532_ hold1929/X _17631_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10744_ hold5725/X _11222_/B _10743_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _10744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _17432_/CLK _16251_/D vssd1 vssd1 vccd1 vccd1 _16251_/Q sky130_fd_sc_hd__dfxtp_1
X_13463_ hold2034/X hold4975/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10675_ hold5617/X _09992_/B _10674_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10675_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ hold1408/X _15221_/B _15201_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _15202_/X
+ sky130_fd_sc_hd__o211a_1
X_12414_ _12426_/A _12414_/B vssd1 vssd1 vccd1 vccd1 _17300_/D sky130_fd_sc_hd__and2_1
X_16182_ _17484_/CLK _16182_/D vssd1 vssd1 vccd1 vccd1 _16182_/Q sky130_fd_sc_hd__dfxtp_1
X_13394_ hold810/X hold4041/X _13844_/C vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _15187_/A _15149_/B vssd1 vssd1 vccd1 vccd1 _15133_/X sky130_fd_sc_hd__or2_1
X_12345_ hold3796/X _12279_/A _12344_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ _15064_/A _15064_/B vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__and2_1
X_12276_ _12282_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ hold2658/X _14040_/B _14014_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14015_/X
+ sky130_fd_sc_hd__o211a_1
X_11227_ _12343_/A _11227_/B vssd1 vssd1 vccd1 vccd1 _11227_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _11203_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _11158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ hold1438/X hold3693/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__mux2_1
X_15966_ _17289_/CLK _15966_/D vssd1 vssd1 vccd1 vccd1 hold549/A sky130_fd_sc_hd__dfxtp_1
X_11089_ hold5431/X _11216_/B _11088_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o211a_1
X_14917_ hold1379/X _14952_/B _14916_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _14917_/X
+ sky130_fd_sc_hd__o211a_1
X_17705_ _17737_/CLK _17705_/D vssd1 vssd1 vccd1 vccd1 _17705_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _17343_/CLK _15897_/D vssd1 vssd1 vccd1 vccd1 hold434/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14848_ _15187_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17636_ _17669_/CLK _17636_/D vssd1 vssd1 vccd1 vccd1 _17636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _17697_/CLK _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
X_14779_ hold1495/X _14772_/B _14778_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14779_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _18080_/CLK _16518_/D vssd1 vssd1 vccd1 vccd1 _16518_/Q sky130_fd_sc_hd__dfxtp_1
X_17498_ _18013_/CLK _17498_/D vssd1 vssd1 vccd1 vccd1 _17498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16449_ _18330_/CLK _16449_/D vssd1 vssd1 vccd1 vccd1 _16449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18119_ _18268_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5605 _11275_/X vssd1 vssd1 vccd1 vccd1 _16915_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5616 _09832_/X vssd1 vssd1 vccd1 vccd1 _16434_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5627 _16891_/Q vssd1 vssd1 vccd1 vccd1 hold5627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5638 _12037_/X vssd1 vssd1 vccd1 vccd1 _17169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4904 _12232_/X vssd1 vssd1 vccd1 vccd1 _17234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5649 _16877_/Q vssd1 vssd1 vccd1 vccd1 hold5649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4915 _17145_/Q vssd1 vssd1 vccd1 vccd1 hold4915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4926 _12286_/X vssd1 vssd1 vccd1 vccd1 _17252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4937 _17281_/Q vssd1 vssd1 vccd1 vccd1 hold4937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4948 _11335_/X vssd1 vssd1 vccd1 vccd1 _16935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4959 _17692_/Q vssd1 vssd1 vccd1 vccd1 hold4959/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout404 hold274/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__buf_6
Xfanout415 _14138_/B vssd1 vssd1 vccd1 vccd1 _14160_/B sky130_fd_sc_hd__buf_6
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout426 _13946_/Y vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__clkbuf_8
X_09823_ hold5419/X _10013_/B _09822_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09823_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout437 fanout484/X vssd1 vssd1 vccd1 vccd1 _13808_/C sky130_fd_sc_hd__buf_4
Xfanout448 _11717_/C vssd1 vssd1 vccd1 vccd1 _12305_/C sky130_fd_sc_hd__clkbuf_8
Xfanout459 _13847_/C vssd1 vssd1 vccd1 vccd1 _13868_/C sky130_fd_sc_hd__clkbuf_4
X_09754_ hold4275/X _11177_/B _09753_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_5_20__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_20__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_08705_ hold5/X _15974_/Q _08721_/S vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09685_ hold5187/X _10067_/B _09684_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09685_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _15374_/A _08636_/B vssd1 vssd1 vccd1 vccd1 _15940_/D sky130_fd_sc_hd__and2_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08567_ _12422_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _15907_/D sky130_fd_sc_hd__and2_1
XFILLER_0_162_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08498_ _15123_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ hold1233/X hold3311/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ hold2288/X _09119_/A2 _09118_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09119_/X
+ sky130_fd_sc_hd__o211a_1
X_10391_ hold766/X hold4141/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ hold5021/X _12311_/B _12129_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ hold4917/X _12347_/B _12060_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__o211a_1
Xhold480 input19/X vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ hold2538/X hold3886/X _11210_/C vssd1 vssd1 vccd1 vccd1 _11013_/B sky130_fd_sc_hd__mux2_1
X_15820_ _17669_/CLK hold226/X vssd1 vssd1 vccd1 vccd1 _15820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _17734_/CLK _15751_/D vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12963_ _12987_/A _12963_/B vssd1 vssd1 vccd1 vccd1 _17497_/D sky130_fd_sc_hd__and2_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _09189_/X vssd1 vssd1 vccd1 vccd1 _16206_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 _18122_/Q vssd1 vssd1 vccd1 vccd1 hold1191/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14988_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14702_/X sky130_fd_sc_hd__or2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ hold4856/X _13811_/B _11913_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__o211a_1
X_15682_ _17769_/CLK _15682_/D vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _12918_/A _12894_/B vssd1 vssd1 vccd1 vccd1 _17474_/D sky130_fd_sc_hd__and2_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17428_/CLK _17421_/D vssd1 vssd1 vccd1 vccd1 _17421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ hold2905/X _14666_/B _14632_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _14633_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ hold4569/X _12323_/B _11844_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11845_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17516_/CLK _17352_/D vssd1 vssd1 vccd1 vccd1 _17352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _15492_/A _14573_/B hold1804/X vssd1 vssd1 vccd1 vccd1 _14564_/X sky130_fd_sc_hd__a21o_1
X_11776_ _12343_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__nor2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16303_ _18460_/CLK hold635/X vssd1 vssd1 vccd1 vccd1 _16303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ _13710_/A _13515_/B vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__or2_1
X_17283_ _17283_/CLK _17283_/D vssd1 vssd1 vccd1 vccd1 _17283_/Q sky130_fd_sc_hd__dfxtp_1
X_10727_ hold886/X _16733_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__mux2_1
X_14495_ hold799/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14495_/X sky130_fd_sc_hd__or2_1
X_16234_ _17754_/CLK _16234_/D vssd1 vssd1 vccd1 vccd1 _16234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13446_ _13734_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10658_ hold1979/X _16710_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _18013_/CLK _16165_/D vssd1 vssd1 vccd1 vccd1 _16165_/Q sky130_fd_sc_hd__dfxtp_1
X_13377_ _13764_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _13377_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _16687_/Q _10589_/B _10589_/C vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__and3_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15116_ hold2058/X _15113_/B _15115_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15116_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ _13873_/A _12328_/B vssd1 vssd1 vccd1 vccd1 _12328_/Y sky130_fd_sc_hd__nor2_1
X_16096_ _16096_/CLK _16096_/D vssd1 vssd1 vccd1 vccd1 hold304/A sky130_fd_sc_hd__dfxtp_1
X_15047_ _15535_/A hold1670/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15048_/B sky130_fd_sc_hd__mux2_1
X_12259_ hold4973/X _12314_/B _12258_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _12259_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2809 _17924_/Q vssd1 vssd1 vccd1 vccd1 hold2809/X sky130_fd_sc_hd__dlygate4sd3_1
X_16998_ _17878_/CLK _16998_/D vssd1 vssd1 vccd1 vccd1 _16998_/Q sky130_fd_sc_hd__dfxtp_1
X_15949_ _17318_/CLK _15949_/D vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ _09471_/B _09481_/B _09470_/C vssd1 vssd1 vccd1 vccd1 _16317_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08421_ _14529_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17619_ _17737_/CLK _17619_/D vssd1 vssd1 vccd1 vccd1 _17619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08352_ _15521_/A hold2461/X hold122/X vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17496_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08283_ _08504_/A hold207/X vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_5_4__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_4__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
Xhold5402 _09919_/X vssd1 vssd1 vccd1 vccd1 _16463_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5413 _16743_/Q vssd1 vssd1 vccd1 vccd1 hold5413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5424 _10657_/X vssd1 vssd1 vccd1 vccd1 _16709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5435 _16978_/Q vssd1 vssd1 vccd1 vccd1 hold5435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4701 _11431_/X vssd1 vssd1 vccd1 vccd1 _16967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5446 _10768_/X vssd1 vssd1 vccd1 vccd1 _16746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4712 _17179_/Q vssd1 vssd1 vccd1 vccd1 hold4712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5457 _11401_/X vssd1 vssd1 vccd1 vccd1 _16957_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4723 _17239_/Q vssd1 vssd1 vccd1 vccd1 hold4723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5468 _16805_/Q vssd1 vssd1 vccd1 vccd1 hold5468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4734 _12178_/X vssd1 vssd1 vccd1 vccd1 _17216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5479 _11020_/X vssd1 vssd1 vccd1 vccd1 _16830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4745 _17003_/Q vssd1 vssd1 vccd1 vccd1 hold4745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4756 _13747_/X vssd1 vssd1 vccd1 vccd1 _17702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4767 _17028_/Q vssd1 vssd1 vccd1 vccd1 hold4767/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout201 _11210_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4778 _10081_/X vssd1 vssd1 vccd1 vccd1 _16517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout212 _10780_/A2 vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__buf_4
Xhold4789 hold5870/X vssd1 vssd1 vccd1 vccd1 hold5871/A sky130_fd_sc_hd__buf_4
Xfanout223 _10558_/A2 vssd1 vssd1 vccd1 vccd1 _11192_/B sky130_fd_sc_hd__buf_4
Xfanout234 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10465_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout245 _10637_/B vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__buf_4
Xfanout256 _13674_/A vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__clkbuf_2
Xfanout267 _11649_/A vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__clkbuf_4
X_09806_ hold863/X _16426_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__mux2_1
Xfanout278 _12243_/A vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__clkbuf_4
X_07998_ hold1163/X _08033_/B _07997_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07998_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout289 _11115_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__buf_4
X_09737_ hold1893/X _16403_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09668_ hold2232/X _16380_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__mux2_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08619_ hold53/X hold601/X _08619_/S vssd1 vssd1 vccd1 vccd1 hold602/A sky130_fd_sc_hd__mux2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ hold2618/X _16357_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__mux2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ hold969/X _17034_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ hold1169/X _17011_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ hold5318/X _13299_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__mux2_1
X_10512_ _10542_/A _10512_/B vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__or2_1
X_14280_ _14728_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__or2_1
X_11492_ hold1621/X _16988_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ _13311_/A1 _13229_/X _13230_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10443_ _10998_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _17571_/Q _17105_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10374_ _10563_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__or2_1
X_12113_ hold1943/X _17195_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__mux2_1
Xhold5980 _15786_/Q vssd1 vssd1 vccd1 vccd1 hold5980/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5991 data_in[29] vssd1 vssd1 vccd1 vccd1 hold377/A sky130_fd_sc_hd__dlygate4sd3_1
X_17970_ _18190_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
X_13093_ _13092_/X hold3188/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_130_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12044_ hold1405/X _17172_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__mux2_1
X_16921_ _17769_/CLK _16921_/D vssd1 vssd1 vccd1 vccd1 _16921_/Q sky130_fd_sc_hd__dfxtp_1
X_16852_ _18055_/CLK _16852_/D vssd1 vssd1 vccd1 vccd1 _16852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout790 fanout842/X vssd1 vssd1 vccd1 vccd1 _08257_/C1 sky130_fd_sc_hd__buf_4
X_15803_ _17747_/CLK _15803_/D vssd1 vssd1 vccd1 vccd1 hold910/A sky130_fd_sc_hd__dfxtp_1
X_16783_ _18062_/CLK _16783_/D vssd1 vssd1 vccd1 vccd1 _16783_/Q sky130_fd_sc_hd__dfxtp_1
X_13995_ hold2328/X _13986_/B _13994_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _13995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15734_ _17737_/CLK _15734_/D vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ hold1237/X _17493_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__mux2_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _17592_/CLK _15665_/D vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfxtp_1
X_18453_ _18454_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
X_12877_ hold1907/X hold3246/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__mux2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _15225_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14616_/X sky130_fd_sc_hd__or2_1
X_17404_ _18456_/CLK _17404_/D vssd1 vssd1 vccd1 vccd1 _17404_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _18390_/CLK hold840/X vssd1 vssd1 vccd1 vccd1 hold839/A sky130_fd_sc_hd__dfxtp_1
X_11828_ hold919/X hold3141/X _12308_/C vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__mux2_1
X_15596_ _17584_/CLK _15596_/D vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17523_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _17335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ _14726_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__or2_1
X_11759_ _11759_/A _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__and3_1
XFILLER_0_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _17266_/CLK _17266_/D vssd1 vssd1 vccd1 vccd1 _17266_/Q sky130_fd_sc_hd__dfxtp_1
X_14478_ hold5971/X _14481_/B _14477_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 hold790/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16217_ _17692_/CLK _16217_/D vssd1 vssd1 vccd1 vccd1 _16217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13429_ hold4893/X _13808_/B _13428_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17197_ _17252_/CLK _17197_/D vssd1 vssd1 vccd1 vccd1 _17197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16148_ _17300_/CLK _16148_/D vssd1 vssd1 vccd1 vccd1 hold397/A sky130_fd_sc_hd__dfxtp_1
Xhold4008 _16985_/Q vssd1 vssd1 vccd1 vccd1 hold4008/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_171_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4019 _10324_/X vssd1 vssd1 vccd1 vccd1 _16598_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _16102_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_100_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18414_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _18410_/CLK _16079_/D vssd1 vssd1 vccd1 vccd1 hold496/A sky130_fd_sc_hd__dfxtp_1
Xhold3307 _16434_/Q vssd1 vssd1 vccd1 vccd1 hold3307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3318 _17282_/Q vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3329 _09676_/X vssd1 vssd1 vccd1 vccd1 _16382_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2606 _09197_/X vssd1 vssd1 vccd1 vccd1 _16210_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07921_ hold1834/X _07924_/B _07920_/Y _08109_/A vssd1 vssd1 vccd1 vccd1 _07921_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2617 _14027_/X vssd1 vssd1 vccd1 vccd1 _17819_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 _16151_/Q vssd1 vssd1 vccd1 vccd1 hold2628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2639 _15747_/Q vssd1 vssd1 vccd1 vccd1 hold2639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 _18129_/Q vssd1 vssd1 vccd1 vccd1 hold1905/X sky130_fd_sc_hd__dlygate4sd3_1
X_07852_ hold1948/X _07869_/B _07851_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _07852_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1916 _07808_/X vssd1 vssd1 vccd1 vccd1 _17752_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1927 _18239_/Q vssd1 vssd1 vccd1 vccd1 hold1927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1938 _17990_/Q vssd1 vssd1 vccd1 vccd1 hold1938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1949 _07852_/X vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 input1/A vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_07783_ hold265/X vssd1 vssd1 vccd1 vccd1 _07783_/Y sky130_fd_sc_hd__inv_2
X_09522_ _09948_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__or2_1
X_09453_ _09456_/B _09456_/C _09456_/D vssd1 vssd1 vccd1 vccd1 _09455_/B sky130_fd_sc_hd__and3_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ hold1366/X _08440_/A2 _08403_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _08404_/X
+ sky130_fd_sc_hd__o211a_1
X_09384_ hold513/X _15474_/B _09383_/X _18460_/Q vssd1 vssd1 vccd1 vccd1 _09384_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _14786_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ _15545_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_259_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17728_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08197_ _14866_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08197_/X sky130_fd_sc_hd__or2_1
Xhold5210 _13789_/X vssd1 vssd1 vccd1 vccd1 _17716_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5221 _16335_/Q vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5232 _10009_/Y vssd1 vssd1 vccd1 vccd1 _16493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5243 _10020_/Y vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5254 _16722_/Q vssd1 vssd1 vccd1 vccd1 hold5254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4520 _17687_/Q vssd1 vssd1 vccd1 vccd1 hold4520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5265 _11197_/Y vssd1 vssd1 vccd1 vccd1 _16889_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4531 _12271_/X vssd1 vssd1 vccd1 vccd1 _17247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5276 _09999_/Y vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5287 _16327_/Q vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__buf_1
Xhold4542 _16566_/Q vssd1 vssd1 vccd1 vccd1 hold4542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4553 _17187_/Q vssd1 vssd1 vccd1 vccd1 hold4553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5298 _11199_/Y vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4564 _13531_/X vssd1 vssd1 vccd1 vccd1 _17630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4575 _16698_/Q vssd1 vssd1 vccd1 vccd1 hold4575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3830 _12373_/Y vssd1 vssd1 vccd1 vccd1 _17281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3841 _16930_/Q vssd1 vssd1 vccd1 vccd1 hold3841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4586 _11299_/X vssd1 vssd1 vccd1 vccd1 _16923_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10090_ hold4830/X _10568_/B _10089_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _16520_/D
+ sky130_fd_sc_hd__o211a_1
Xhold3852 _16525_/Q vssd1 vssd1 vccd1 vccd1 hold3852/X sky130_fd_sc_hd__clkbuf_2
Xhold4597 _17148_/Q vssd1 vssd1 vccd1 vccd1 hold4597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3863 _16427_/Q vssd1 vssd1 vccd1 vccd1 hold3863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3874 hold4679/X vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3885 _13813_/Y vssd1 vssd1 vccd1 vccd1 _17724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3896 _13837_/Y vssd1 vssd1 vccd1 vccd1 _17732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ hold3087/X _12799_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__mux2_1
X_13780_ _13874_/A _13886_/B _13779_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13780_/X
+ sky130_fd_sc_hd__o211a_1
X_10992_ _11121_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ hold3468/X _12730_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ hold631/X _15485_/A2 _15485_/B1 hold700/X _15448_/X vssd1 vssd1 vccd1 vccd1
+ _15452_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ hold3103/X _12661_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__mux2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _15189_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14401_/X sky130_fd_sc_hd__or2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _12093_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__or2_1
X_15381_ _16302_/Q _09362_/A _09392_/B hold535/X _15380_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_53_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12593_ hold3435/X _12592_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17120_ _17283_/CLK _17120_/D vssd1 vssd1 vccd1 vccd1 _17120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14332_ _14726_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11544_ _11640_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17051_ _17908_/CLK _17051_/D vssd1 vssd1 vccd1 vccd1 _17051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ hold2308/X _14272_/B _14262_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _14263_/X
+ sky130_fd_sc_hd__o211a_1
X_11475_ _11667_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__or2_1
X_16002_ _18409_/CLK _16002_/D vssd1 vssd1 vccd1 vccd1 _16002_/Q sky130_fd_sc_hd__dfxtp_1
X_13214_ _13214_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13214_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ hold3924/X _10897_/A2 _10425_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _10426_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ hold466/X _14214_/B vssd1 vssd1 vccd1 vccd1 hold467/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _13145_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10357_ hold4016/X _10643_/B _10356_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ hold4987/X _13075_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17953_ _18391_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
X_10288_ hold3558/X _10558_/A2 _10287_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10288_/X
+ sky130_fd_sc_hd__o211a_1
X_12027_ _12285_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__or2_1
X_16904_ _17879_/CLK _16904_/D vssd1 vssd1 vccd1 vccd1 _16904_/Q sky130_fd_sc_hd__dfxtp_1
X_17884_ _17884_/CLK hold872/X vssd1 vssd1 vccd1 vccd1 hold871/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ _18070_/CLK _16835_/D vssd1 vssd1 vccd1 vccd1 _16835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _15105_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__or2_1
X_16766_ _18025_/CLK _16766_/D vssd1 vssd1 vccd1 vccd1 _16766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15717_ _17253_/CLK _15717_/D vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfxtp_1
X_12929_ hold3584/X _12928_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__mux2_1
X_16697_ _18095_/CLK _16697_/D vssd1 vssd1 vccd1 vccd1 _16697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18436_ _18441_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
X_15648_ _17128_/CLK _15648_/D vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15579_ _17282_/CLK _15579_/D vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfxtp_1
X_18367_ _18391_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ _15525_/A hold2468/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__mux2_1
X_17318_ _17318_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 _17318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _18330_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08051_ hold2397/X _08082_/B _08050_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08051_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17249_ _17281_/CLK _17249_/D vssd1 vssd1 vccd1 vccd1 _17249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3104 _17496_/Q vssd1 vssd1 vccd1 vccd1 hold3104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3115 hold5852/X vssd1 vssd1 vccd1 vccd1 hold5853/A sky130_fd_sc_hd__buf_4
Xhold3126 _16547_/Q vssd1 vssd1 vccd1 vccd1 hold3126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ hold443/X hold495/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__mux2_1
Xhold3137 _10612_/Y vssd1 vssd1 vccd1 vccd1 _16694_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3148 _12369_/Y vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2403 _18100_/Q vssd1 vssd1 vccd1 vccd1 hold2403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3159 _17568_/Q vssd1 vssd1 vccd1 vccd1 hold3159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 _12590_/X vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _15844_/Q vssd1 vssd1 vccd1 vccd1 hold2425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2436 _08461_/X vssd1 vssd1 vccd1 vccd1 _15859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07904_ _15527_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1702 _18235_/Q vssd1 vssd1 vccd1 vccd1 hold1702/X sky130_fd_sc_hd__dlygate4sd3_1
X_08884_ hold47/X hold567/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__mux2_1
Xhold2447 _16259_/Q vssd1 vssd1 vccd1 vccd1 hold2447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1713 _07913_/X vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 _09143_/X vssd1 vssd1 vccd1 vccd1 _16184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 _14637_/X vssd1 vssd1 vccd1 vccd1 _18111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2469 _15684_/Q vssd1 vssd1 vccd1 vccd1 hold2469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1735 _14137_/X vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1746 _18214_/Q vssd1 vssd1 vccd1 vccd1 hold1746/X sky130_fd_sc_hd__dlygate4sd3_1
X_07835_ _14740_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07835_/X sky130_fd_sc_hd__or2_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1757 _09429_/X vssd1 vssd1 vccd1 vccd1 _16300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1768 _18387_/Q vssd1 vssd1 vccd1 vccd1 hold1768/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 _14422_/X vssd1 vssd1 vccd1 vccd1 _18009_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09505_ hold5532/X _09998_/B _09504_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _09505_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ hold616/X _16304_/Q vssd1 vssd1 vccd1 vccd1 hold617/A sky130_fd_sc_hd__or2_1
XFILLER_0_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A _09386_/D vssd1 vssd1 vccd1 vccd1 _09369_/D sky130_fd_sc_hd__or2_1
XFILLER_0_118_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ hold2028/X _08323_/B _08317_/Y _12756_/A vssd1 vssd1 vccd1 vccd1 _08318_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 _15515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ hold2447/X _09338_/A2 _09297_/X _12927_/A vssd1 vssd1 vccd1 vccd1 _09298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_61 hold173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_72 hold800/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08249_ hold2637/X _08268_/B _08248_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08249_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_83 hold5853/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_94 _14286_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ hold4020/X _11747_/B _11259_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5040 _16379_/Q vssd1 vssd1 vccd1 vccd1 hold5040/X sky130_fd_sc_hd__dlygate4sd3_1
X_10211_ hold2203/X hold4407/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__mux2_1
Xhold5051 _11005_/X vssd1 vssd1 vccd1 vccd1 _16825_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5062 _17737_/Q vssd1 vssd1 vccd1 vccd1 hold5062/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5073 _09856_/X vssd1 vssd1 vccd1 vccd1 _16442_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11191_ _11218_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11191_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5084 _16755_/Q vssd1 vssd1 vccd1 vccd1 hold5084/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4350 _10111_/X vssd1 vssd1 vccd1 vccd1 _16527_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5095 _10087_/X vssd1 vssd1 vccd1 vccd1 _16519_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4361 _16672_/Q vssd1 vssd1 vccd1 vccd1 hold4361/X sky130_fd_sc_hd__dlygate4sd3_1
X_10142_ hold1161/X hold3745/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__mux2_1
Xhold4372 _10762_/X vssd1 vssd1 vccd1 vccd1 _16744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4383 _17629_/Q vssd1 vssd1 vccd1 vccd1 hold4383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4394 _12112_/X vssd1 vssd1 vccd1 vccd1 _17194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3660 _10053_/Y vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14950_ _14950_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14950_/Y sky130_fd_sc_hd__nand2_1
X_10073_ _16515_/Q _10073_/B _10481_/S vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__and3_1
Xhold3671 _13830_/Y vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3682 _10041_/Y vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3693 _16527_/Q vssd1 vssd1 vccd1 vccd1 hold3693/X sky130_fd_sc_hd__buf_2
X_13901_ _13901_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _17758_/D sky130_fd_sc_hd__and2_1
Xhold2970 _14552_/X vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14881_ hold2445/X _14880_/B _14880_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14881_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2981 _18353_/Q vssd1 vssd1 vccd1 vccd1 hold2981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2992 _18053_/Q vssd1 vssd1 vccd1 vccd1 hold2992/X sky130_fd_sc_hd__dlygate4sd3_1
X_16620_ _18210_/CLK _16620_/D vssd1 vssd1 vccd1 vccd1 _16620_/Q sky130_fd_sc_hd__dfxtp_1
X_13832_ _17731_/Q _13832_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16551_ _18205_/CLK _16551_/D vssd1 vssd1 vccd1 vccd1 _16551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13763_ hold1765/X hold5156/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13764_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ hold5741/X _11201_/B _10974_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _10975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _12777_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _17414_/D sky130_fd_sc_hd__and2_1
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__and2_1
X_16482_ _18395_/CLK _16482_/D vssd1 vssd1 vccd1 vccd1 _16482_/Q sky130_fd_sc_hd__dfxtp_1
X_13694_ hold2008/X hold3513/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18221_ _18221_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_15433_ _15481_/A1 _15425_/X _15432_/X _15481_/B1 _18419_/Q vssd1 vssd1 vccd1 vccd1
+ _15433_/X sky130_fd_sc_hd__a32o_1
X_12645_ _12876_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__and2_1
XFILLER_0_155_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15364_ _15364_/A _15364_/B vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__and2_1
X_18152_ _18216_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_12576_ _12987_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _17368_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17103_ _17276_/CLK _17103_/D vssd1 vssd1 vccd1 vccd1 _17103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14315_ hold1665/X _14333_/A2 _14314_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _14315_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18083_ _18266_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
X_11527_ hold4860/X _12299_/B _11526_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11527_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ hold706/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17034_ _17882_/CLK _17034_/D vssd1 vssd1 vccd1 vccd1 _17034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14246_ _14246_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ hold4469/X _12320_/B _11457_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10409_ hold2274/X hold4435/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177_ hold2783/X _14198_/B _14176_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14177_/X
+ sky130_fd_sc_hd__o211a_1
X_11389_ hold4008/X _12338_/B _11388_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 _11389_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13121_/X _13127_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17534_/D sky130_fd_sc_hd__o21a_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13058_/X _16900_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
X_17936_ _18025_/CLK hold887/X vssd1 vssd1 vccd1 vccd1 hold886/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1009 _07840_/X vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17867_ _17908_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16818_ _18053_/CLK _16818_/D vssd1 vssd1 vccd1 vccd1 _16818_/Q sky130_fd_sc_hd__dfxtp_1
X_17798_ _17798_/CLK hold976/X vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16749_ _17984_/CLK _16749_/D vssd1 vssd1 vccd1 vccd1 _16749_/Q sky130_fd_sc_hd__dfxtp_1
X_09221_ hold1994/X _09216_/B _09220_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _09221_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18419_ _18423_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _15535_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08103_ hold816/A hold281/A vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ hold1237/X _09119_/A2 _09082_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _09083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08034_ hold2239/X _08033_/B _08033_/Y _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08034_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput70 input70/A vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 hold832/A vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold843 hold843/A vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 hold854/A vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/A vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/A vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold887 hold887/A vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 input3/X vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _13070_/A _10016_/B _09984_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _16485_/D
+ sky130_fd_sc_hd__o211a_1
Xhold2200 _08330_/X vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2211 input69/X vssd1 vssd1 vccd1 vccd1 hold2211/X sky130_fd_sc_hd__dlygate4sd3_1
X_08936_ _13002_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _16085_/D sky130_fd_sc_hd__and2_1
Xhold2222 _15657_/Q vssd1 vssd1 vccd1 vccd1 hold2222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2233 _15015_/X vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2244 _18458_/Q vssd1 vssd1 vccd1 vccd1 hold2244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 _07882_/X vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 _08273_/X vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _17945_/Q vssd1 vssd1 vccd1 vccd1 hold1521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2266 _18210_/Q vssd1 vssd1 vccd1 vccd1 hold2266/X sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ _09063_/A hold566/X vssd1 vssd1 vccd1 vccd1 _16052_/D sky130_fd_sc_hd__and2_1
Xhold1532 _14859_/X vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 _18116_/Q vssd1 vssd1 vccd1 vccd1 hold2277/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1543 _14303_/X vssd1 vssd1 vccd1 vccd1 _17951_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2288 _16174_/Q vssd1 vssd1 vccd1 vccd1 hold2288/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2299 _14329_/X vssd1 vssd1 vccd1 vccd1 _17964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _14319_/X vssd1 vssd1 vccd1 vccd1 _17959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 _18191_/Q vssd1 vssd1 vccd1 vccd1 hold1565/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1576 _18238_/Q vssd1 vssd1 vccd1 vccd1 hold1576/X sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ hold624/A hold606/A hold298/A hold279/X vssd1 vssd1 vccd1 vccd1 _14735_/A
+ sky130_fd_sc_hd__or4bb_4
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _15491_/A hold705/X vssd1 vssd1 vccd1 vccd1 _16018_/D sky130_fd_sc_hd__and2_1
Xhold1587 _18326_/Q vssd1 vssd1 vccd1 vccd1 hold1587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1598 _14589_/X vssd1 vssd1 vccd1 vccd1 _18088_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ hold689/X _16744_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_274_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ _07804_/A _09463_/C _15304_/A _09418_/X vssd1 vssd1 vccd1 vccd1 _09419_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_203_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10691_ hold2809/X hold3129/X _11210_/C vssd1 vssd1 vccd1 vccd1 _10692_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _17308_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _13873_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14100_ _15553_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14100_/X sky130_fd_sc_hd__or2_1
X_11312_ hold1334/X hold3713/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__mux2_1
X_15080_ hold1523/X _15113_/B _15079_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15080_/X
+ sky130_fd_sc_hd__o211a_1
X_12292_ hold4447/X _12308_/B _12291_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o211a_1
X_14031_ hold2147/X _14036_/B _14030_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14031_/X
+ sky130_fd_sc_hd__o211a_1
X_11243_ _18431_/Q hold3787/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__mux2_1
X_11174_ _16882_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__and3_1
Xhold4180 _16692_/Q vssd1 vssd1 vccd1 vccd1 hold4180/X sky130_fd_sc_hd__dlygate4sd3_1
X_10125_ _10551_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__or2_1
Xhold4191 _10102_/X vssd1 vssd1 vccd1 vccd1 _16524_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15982_ _17307_/CLK _15982_/D vssd1 vssd1 vccd1 vccd1 hold450/A sky130_fd_sc_hd__dfxtp_1
Xhold3490 _12719_/X vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17721_ _17721_/CLK _17721_/D vssd1 vssd1 vccd1 vccd1 _17721_/Q sky130_fd_sc_hd__dfxtp_1
X_10056_ _13262_/A _09954_/A _10055_/X vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__a21oi_1
X_14933_ hold1220/X _14952_/B _14932_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17652_ _17748_/CLK _17652_/D vssd1 vssd1 vccd1 vccd1 _17652_/Q sky130_fd_sc_hd__dfxtp_1
X_14864_ _14988_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__or2_1
X_16603_ _18225_/CLK _16603_/D vssd1 vssd1 vccd1 vccd1 _16603_/Q sky130_fd_sc_hd__dfxtp_1
X_13815_ hold3622/X _13713_/A _13814_/X vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__a21oi_1
X_14795_ hold5957/X _14822_/B hold1059/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14795_/X
+ sky130_fd_sc_hd__o211a_1
X_17583_ _17583_/CLK _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13746_ _13764_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__or2_1
X_16534_ _18140_/CLK _16534_/D vssd1 vssd1 vccd1 vccd1 _16534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ hold1925/X _16810_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _18378_/CLK _16465_/D vssd1 vssd1 vccd1 vccd1 _16465_/Q sky130_fd_sc_hd__dfxtp_1
X_13677_ _13776_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10889_ hold1938/X _16787_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18204_ _18204_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
X_15416_ _17317_/Q _15479_/A2 _09392_/A hold696/X vssd1 vssd1 vccd1 vccd1 _15416_/X
+ sky130_fd_sc_hd__a22o_1
X_12628_ hold2557/X hold3072/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12628_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16396_ _18334_/CLK _16396_/D vssd1 vssd1 vccd1 vccd1 _16396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ hold477/X _15479_/A2 _09386_/D hold640/X _15346_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18135_ _18231_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12559_ hold2701/X _17364_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5809 output96/X vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15278_ hold238/X _15484_/A2 _15451_/A2 hold449/X vssd1 vssd1 vccd1 vccd1 _15278_/X
+ sky130_fd_sc_hd__a22o_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
X_18066_ _18066_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold478/X vssd1 vssd1 vccd1 vccd1 hold479/A sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _17769_/CLK _17017_/D vssd1 vssd1 vccd1 vccd1 _17017_/Q sky130_fd_sc_hd__dfxtp_1
X_14229_ hold1018/X _14216_/Y _14228_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14229_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_78_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17525_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout608 _15447_/B1 vssd1 vssd1 vccd1 vccd1 _09392_/C sky130_fd_sc_hd__buf_6
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _09354_/Y vssd1 vssd1 vccd1 vccd1 _15479_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ hold2926/X hold3328/X _11177_/C vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__mux2_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ hold359/X hold450/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__mux2_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _18273_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_1
X_08652_ _15354_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _15948_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08583_ _15304_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _15915_/D sky130_fd_sc_hd__and2_1
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09204_ _15533_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ hold1263/X _09177_/A2 _09134_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _15182_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _09066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ _15531_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__or2_1
Xhold640 hold640/A vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold651 hold651/A vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 hold673/A vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 hold684/A vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 hold695/A vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09968_ hold930/X _16480_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__mux2_1
Xhold2030 _16273_/Q vssd1 vssd1 vccd1 vccd1 hold2030/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2041 _08071_/X vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _12430_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _16077_/D sky130_fd_sc_hd__and2_1
Xhold2052 _18016_/Q vssd1 vssd1 vccd1 vccd1 hold2052/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2063 _15546_/X vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 _18286_/Q vssd1 vssd1 vccd1 vccd1 hold2074/X sky130_fd_sc_hd__dlygate4sd3_1
X_09899_ hold853/X _16457_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__mux2_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2085 _15742_/Q vssd1 vssd1 vccd1 vccd1 hold2085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1340 hold1340/A vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ hold2574/X _17134_/Q _12353_/C vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__mux2_1
Xhold1351 _17842_/Q vssd1 vssd1 vccd1 vccd1 hold1351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2096 _17969_/Q vssd1 vssd1 vccd1 vccd1 hold2096/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 _09195_/X vssd1 vssd1 vccd1 vccd1 _16209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 _18268_/Q vssd1 vssd1 vccd1 vccd1 hold1373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 _14025_/X vssd1 vssd1 vccd1 vccd1 _17818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1395 _15639_/Q vssd1 vssd1 vccd1 vccd1 hold1395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ hold2480/X hold3877/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ hold3513/X _13880_/B _13599_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13600_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _11097_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__or2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14580_ _15189_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11792_ _17088_/Q _11792_/B _11792_/C vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__and3_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ hold4563/X _13829_/B _13530_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10743_ _11694_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _17447_/CLK _16250_/D vssd1 vssd1 vccd1 vccd1 _16250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13462_ hold3577/X _13886_/B _13461_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13462_/X
+ sky130_fd_sc_hd__o211a_1
X_10674_ _11067_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10674_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15201_ hold883/X _15233_/B vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__or2_1
X_12413_ hold214/X hold395/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__mux2_1
X_16181_ _17464_/CLK _16181_/D vssd1 vssd1 vccd1 vccd1 _16181_/Q sky130_fd_sc_hd__dfxtp_1
X_13393_ hold4589/X _13856_/B _13392_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15132_ hold1589/X _15161_/B _15131_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _15132_/X
+ sky130_fd_sc_hd__o211a_1
X_12344_ _17272_/Q _13844_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15063_ _15225_/A hold1477/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15064_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12275_ hold1960/X hold4536/X _12377_/C vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__mux2_1
X_14014_ _15521_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14014_/X sky130_fd_sc_hd__or2_1
X_11226_ hold5300/X _11670_/A _11225_/X vssd1 vssd1 vccd1 vccd1 _11226_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ hold3636/X _11136_/A _11156_/X vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10108_ hold4891/X _10628_/B _10107_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__o211a_1
X_15965_ _17284_/CLK _15965_/D vssd1 vssd1 vccd1 vccd1 hold426/A sky130_fd_sc_hd__dfxtp_1
X_11088_ _11121_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__or2_1
X_17704_ _17738_/CLK _17704_/D vssd1 vssd1 vccd1 vccd1 _17704_/Q sky130_fd_sc_hd__dfxtp_1
X_10039_ _10588_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _16503_/D sky130_fd_sc_hd__nor2_1
X_14916_ _14970_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14916_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_196_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18020_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15896_ _17314_/CLK _15896_/D vssd1 vssd1 vccd1 vccd1 hold519/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _17669_/CLK _17635_/D vssd1 vssd1 vccd1 vccd1 _17635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ hold1499/X _14880_/B _14846_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_125_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18395_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _17686_/CLK _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
X_14778_ _15225_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16517_ _18267_/CLK _16517_/D vssd1 vssd1 vccd1 vccd1 _16517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ hold4682/X _13832_/B _13728_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13729_/X
+ sky130_fd_sc_hd__o211a_1
X_17497_ _17981_/CLK _17497_/D vssd1 vssd1 vccd1 vccd1 _17497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ _18235_/CLK _16448_/D vssd1 vssd1 vccd1 vccd1 _16448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_5_3__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16379_ _18355_/CLK _16379_/D vssd1 vssd1 vccd1 vccd1 _16379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18118_ _18118_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5606 _16875_/Q vssd1 vssd1 vccd1 vccd1 hold5606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5617 _16747_/Q vssd1 vssd1 vccd1 vccd1 hold5617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5628 _11107_/X vssd1 vssd1 vccd1 vccd1 _16859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5639 _16370_/Q vssd1 vssd1 vccd1 vccd1 hold5639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4905 _17224_/Q vssd1 vssd1 vccd1 vccd1 hold4905/X sky130_fd_sc_hd__dlygate4sd3_1
X_18049_ _18050_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4916 _11869_/X vssd1 vssd1 vccd1 vccd1 _17113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4927 _17063_/Q vssd1 vssd1 vccd1 vccd1 hold4927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4938 _12277_/X vssd1 vssd1 vccd1 vccd1 _17249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4949 _17749_/Q vssd1 vssd1 vccd1 vccd1 hold4949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout405 hold274/X vssd1 vssd1 vccd1 vccd1 _14391_/S sky130_fd_sc_hd__clkbuf_8
Xfanout416 hold586/X vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__clkbuf_8
X_09822_ _09918_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__or2_1
Xfanout427 hold243/X vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__buf_6
Xfanout438 _12308_/C vssd1 vssd1 vccd1 vccd1 _13811_/C sky130_fd_sc_hd__clkbuf_8
Xfanout449 _11717_/C vssd1 vssd1 vccd1 vccd1 _11732_/C sky130_fd_sc_hd__clkbuf_8
X_09753_ _11082_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09753_/X sky130_fd_sc_hd__or2_1
X_08704_ _12438_/A _08704_/B vssd1 vssd1 vccd1 vccd1 _15973_/D sky130_fd_sc_hd__and2_1
XFILLER_0_193_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09684_ _10491_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ hold219/X hold721/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08636_/B sky130_fd_sc_hd__mux2_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ hold184/X hold651/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__mux2_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08497_ hold2555/X _08486_/B _08496_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08497_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09118_ _15559_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10390_ hold4079/X _10580_/B _10389_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09049_ _15334_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _16141_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12060_ _12255_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__or2_1
Xhold470 hold470/A vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ hold5554/X _11201_/B _11010_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o211a_1
Xhold492 hold492/A vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _17669_/CLK _15750_/D vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfxtp_1
X_12962_ hold3084/X _12961_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__mux2_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _14111_/X vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _18252_/Q vssd1 vssd1 vccd1 vccd1 hold1181/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ hold2907/X _14720_/B _14700_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _14701_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _13716_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__or2_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1192 _14659_/X vssd1 vssd1 vccd1 vccd1 _18122_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _17905_/CLK _15681_/D vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfxtp_1
X_12893_ hold3018/X _12892_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__mux2_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17428_/CLK _17420_/D vssd1 vssd1 vccd1 vccd1 _17420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14740_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__or2_1
X_11844_ _12036_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17513_/CLK _17351_/D vssd1 vssd1 vccd1 vccd1 _17351_/Q sky130_fd_sc_hd__dfxtp_1
X_14563_ _14740_/A _14557_/Y hold1795/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _14563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11775_ hold5289/X _12051_/A _11774_/X vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__a21oi_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _18460_/CLK hold630/X vssd1 vssd1 vccd1 vccd1 _16302_/Q sky130_fd_sc_hd__dfxtp_1
X_13514_ hold2561/X hold4836/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__mux2_1
X_10726_ hold5546/X _11762_/B _10725_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _10726_/X
+ sky130_fd_sc_hd__o211a_1
X_17282_ _17282_/CLK _17282_/D vssd1 vssd1 vccd1 vccd1 _17282_/Q sky130_fd_sc_hd__dfxtp_1
X_14494_ hold954/X _14487_/B _14493_/X _14362_/A vssd1 vssd1 vccd1 vccd1 hold955/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16233_ _17435_/CLK _16233_/D vssd1 vssd1 vccd1 vccd1 _16233_/Q sky130_fd_sc_hd__dfxtp_1
X_13445_ _15839_/Q _17602_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ hold5423/X _11156_/B _10656_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ hold808/X _17579_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__mux2_1
X_16164_ _18013_/CLK _16164_/D vssd1 vssd1 vccd1 vccd1 _16164_/Q sky130_fd_sc_hd__dfxtp_1
X_10588_ _10588_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ _15169_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15115_/X sky130_fd_sc_hd__or2_1
X_12327_ hold3168/X _12243_/A _12326_/X vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__a21oi_1
X_16095_ _18423_/CLK _16095_/D vssd1 vssd1 vccd1 vccd1 _16095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15046_ _15050_/A _15046_/B vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__and2_1
X_12258_ _13794_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__or2_1
X_11209_ _12343_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11209_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12189_ _13794_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_306_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17693_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16997_ _17877_/CLK _16997_/D vssd1 vssd1 vccd1 vccd1 _16997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _18411_/CLK _15948_/D vssd1 vssd1 vccd1 vccd1 hold554/A sky130_fd_sc_hd__dfxtp_1
X_15879_ _17686_/CLK _15879_/D vssd1 vssd1 vccd1 vccd1 _15879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ hold5951/X _08433_/B hold1099/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08420_/X
+ sky130_fd_sc_hd__o211a_1
X_17618_ _17747_/CLK _17618_/D vssd1 vssd1 vccd1 vccd1 _17618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17549_ _18185_/CLK _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ hold624/A hold606/A hold298/A hold279/X vssd1 vssd1 vccd1 vccd1 hold207/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17375_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5403 _17012_/Q vssd1 vssd1 vccd1 vccd1 hold5403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5414 _10663_/X vssd1 vssd1 vccd1 vccd1 _16711_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5425 _16369_/Q vssd1 vssd1 vccd1 vccd1 hold5425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5436 _11368_/X vssd1 vssd1 vccd1 vccd1 _16946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4702 _17058_/Q vssd1 vssd1 vccd1 vccd1 hold4702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5447 _16733_/Q vssd1 vssd1 vccd1 vccd1 hold5447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5458 _16461_/Q vssd1 vssd1 vccd1 vccd1 hold5458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4713 _11971_/X vssd1 vssd1 vccd1 vccd1 _17147_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4724 _12151_/X vssd1 vssd1 vccd1 vccd1 _17207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5469 _10849_/X vssd1 vssd1 vccd1 vccd1 _16773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4735 _16614_/Q vssd1 vssd1 vccd1 vccd1 hold4735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4746 _11443_/X vssd1 vssd1 vccd1 vccd1 _16971_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4757 _16820_/Q vssd1 vssd1 vccd1 vccd1 hold4757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4768 _11518_/X vssd1 vssd1 vccd1 vccd1 _16996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4779 _16613_/Q vssd1 vssd1 vccd1 vccd1 hold4779/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout202 fanout209/X vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__clkbuf_4
Xfanout213 _10780_/A2 vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__buf_4
Xfanout224 _10465_/A2 vssd1 vssd1 vccd1 vccd1 _10558_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout235 _09952_/A2 vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__buf_4
Xfanout246 _10637_/B vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__buf_4
X_09805_ hold5600/X _09998_/B _09804_/X _14905_/C1 vssd1 vssd1 vccd1 vccd1 _09805_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout257 _13674_/A vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__clkbuf_4
Xfanout268 _11649_/A vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__buf_4
X_07997_ hold756/X _08045_/B vssd1 vssd1 vccd1 vccd1 _07997_/X sky130_fd_sc_hd__or2_1
Xfanout279 fanout298/X vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__clkbuf_4
X_09736_ hold3307/X _10022_/B _09735_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09736_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ hold5009/X _10070_/B _09666_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09667_/X
+ sky130_fd_sc_hd__o211a_1
X_08618_ _09003_/A _08618_/B vssd1 vssd1 vccd1 vccd1 _15931_/D sky130_fd_sc_hd__and2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ hold5695/X _10016_/B _09597_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09598_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _15284_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _15898_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ hold5504/X _12329_/B _11559_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11560_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10511_ hold2736/X hold4057/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ hold4492/X _12320_/B _11490_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11491_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ hold2776/X hold4254/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13161_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__and2_1
X_10373_ hold2730/X hold4883/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12112_ hold4393/X _13811_/B _12111_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _12112_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5970 _17900_/Q vssd1 vssd1 vccd1 vccd1 hold5970/X sky130_fd_sc_hd__dlygate4sd3_1
X_13092_ hold3751/X _13091_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_1
Xhold5981 _16276_/Q vssd1 vssd1 vccd1 vccd1 hold5981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5992 data_in[27] vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dlygate4sd3_1
X_12043_ hold5369/X _12329_/B _12042_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _12043_/X
+ sky130_fd_sc_hd__o211a_1
X_16920_ _17903_/CLK _16920_/D vssd1 vssd1 vccd1 vccd1 _16920_/Q sky130_fd_sc_hd__dfxtp_1
X_16851_ _18054_/CLK _16851_/D vssd1 vssd1 vccd1 vccd1 _16851_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout780 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _14191_/C1 sky130_fd_sc_hd__buf_4
X_15802_ _17735_/CLK _15802_/D vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout791 _15056_/A vssd1 vssd1 vccd1 vccd1 _15168_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16782_ _18337_/CLK _16782_/D vssd1 vssd1 vccd1 vccd1 _16782_/Q sky130_fd_sc_hd__dfxtp_1
X_13994_ _14728_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _17647_/CLK _15733_/D vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _12996_/A _12945_/B vssd1 vssd1 vccd1 vccd1 _17491_/D sky130_fd_sc_hd__and2_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18454_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _17208_/CLK _15664_/D vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12876_/A _12876_/B vssd1 vssd1 vccd1 vccd1 _17468_/D sky130_fd_sc_hd__and2_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _18454_/CLK _17403_/D vssd1 vssd1 vccd1 vccd1 _17403_/Q sky130_fd_sc_hd__dfxtp_1
X_14615_ hold1852/X _14610_/B _14614_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14615_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11827_ hold5028/X _12305_/B _11826_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11827_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18383_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
X_15595_ _17211_/CLK _15595_/D vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17341_/CLK hold220/X vssd1 vssd1 vccd1 vccd1 _17334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11758_ _12331_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11758_/Y sky130_fd_sc_hd__nor2_1
X_14546_ hold1447/X _14541_/B _14545_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ hold2742/X hold5245/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17265_ _17900_/CLK _17265_/D vssd1 vssd1 vccd1 vccd1 _17265_/Q sky130_fd_sc_hd__dfxtp_1
X_11689_ hold4053/X _11783_/B _11688_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11689_/X
+ sky130_fd_sc_hd__o211a_1
X_14477_ hold735/X _14479_/B vssd1 vssd1 vccd1 vccd1 _14477_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16216_ _17692_/CLK _16216_/D vssd1 vssd1 vccd1 vccd1 _16216_/Q sky130_fd_sc_hd__dfxtp_1
X_13428_ _13713_/A _13428_/B vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17196_ _17260_/CLK _17196_/D vssd1 vssd1 vccd1 vccd1 _17196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _17314_/CLK _16147_/D vssd1 vssd1 vccd1 vccd1 hold445/A sky130_fd_sc_hd__dfxtp_1
X_13359_ _13770_/A _13359_/B vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__or2_1
Xhold4009 _11389_/X vssd1 vssd1 vccd1 vccd1 _16953_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3308 _09736_/X vssd1 vssd1 vccd1 vccd1 _16402_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16078_ _17313_/CLK _16078_/D vssd1 vssd1 vccd1 vccd1 hold529/A sky130_fd_sc_hd__dfxtp_1
Xhold3319 _12280_/X vssd1 vssd1 vccd1 vccd1 _17250_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _15543_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07920_/Y sky130_fd_sc_hd__nand2_1
X_15029_ _15191_/A hold1656/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15030_/B sky130_fd_sc_hd__mux2_1
Xhold2607 _17816_/Q vssd1 vssd1 vccd1 vccd1 hold2607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 _18270_/Q vssd1 vssd1 vccd1 vccd1 hold2618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _09073_/X vssd1 vssd1 vccd1 vccd1 _16151_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1906 _14673_/X vssd1 vssd1 vccd1 vccd1 _18129_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07851_ _15529_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07851_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_140_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18396_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1917 _16196_/Q vssd1 vssd1 vccd1 vccd1 hold1917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 _14903_/X vssd1 vssd1 vccd1 vccd1 _18239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _17823_/Q vssd1 vssd1 vccd1 vccd1 hold1939/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput2 input2/A vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_07782_ hold235/X vssd1 vssd1 vccd1 vccd1 _07782_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_190_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ hold2559/X _13118_/A _10001_/C vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09456_/C _09456_/D _09456_/B vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _15517_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09383_ _15489_/A _09383_/B _09383_/C _09383_/D vssd1 vssd1 vccd1 vccd1 _09383_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08334_ hold2553/X _08336_/A2 _08333_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08265_ hold1824/X _08268_/B _08264_/Y _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ hold1891/X _08213_/B _08195_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _08196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5200 _09377_/X vssd1 vssd1 vccd1 vccd1 _16280_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5211 _17747_/Q vssd1 vssd1 vccd1 vccd1 hold5211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5222 _10014_/Y vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5233 _16915_/Q vssd1 vssd1 vccd1 vccd1 hold5233/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_299_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17697_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5244 _10021_/Y vssd1 vssd1 vccd1 vccd1 _16497_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4510 _16659_/Q vssd1 vssd1 vccd1 vccd1 hold4510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5255 _11175_/Y vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4521 _13606_/X vssd1 vssd1 vccd1 vccd1 _17655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5266 _16735_/Q vssd1 vssd1 vccd1 vccd1 hold5266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4532 _17071_/Q vssd1 vssd1 vccd1 vccd1 hold4532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5277 _10000_/Y vssd1 vssd1 vccd1 vccd1 _16490_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5288 _09991_/Y vssd1 vssd1 vccd1 vccd1 _16487_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_228_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17906_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4543 _10132_/X vssd1 vssd1 vccd1 vccd1 _16534_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4554 _11995_/X vssd1 vssd1 vccd1 vccd1 _17155_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3820 _12360_/Y vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5299 _11200_/Y vssd1 vssd1 vccd1 vccd1 _16890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4565 _16651_/Q vssd1 vssd1 vccd1 vccd1 hold4565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3831 _16363_/Q vssd1 vssd1 vccd1 vccd1 hold3831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4576 _10528_/X vssd1 vssd1 vccd1 vccd1 _16666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3842 _11799_/Y vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4587 _16781_/Q vssd1 vssd1 vccd1 vccd1 hold4587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3853 _10584_/Y vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4598 _11878_/X vssd1 vssd1 vccd1 vccd1 _17116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3864 _09715_/X vssd1 vssd1 vccd1 vccd1 _16395_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3875 _10587_/Y vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3886 _16828_/Q vssd1 vssd1 vccd1 vccd1 hold3886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3897 _17116_/Q vssd1 vssd1 vccd1 vccd1 hold3897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ hold1970/X hold3917/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__mux2_1
X_10991_ hold2878/X hold3915/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ hold1575/X hold3085/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__mux2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ hold2357/X hold3055/X _12910_/S vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__mux2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ hold1818/X _17028_/Q _12320_/C vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__mux2_1
X_14400_ hold2760/X hold209/X _14399_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14400_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ hold697/X _09367_/A _09392_/A hold647/X vssd1 vssd1 vccd1 vccd1 _15380_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ hold2030/X hold3375/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ hold1896/X hold4178/X _11735_/C vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__mux2_1
X_14331_ hold1412/X _14326_/B _14330_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14331_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17050_ _17898_/CLK _17050_/D vssd1 vssd1 vccd1 vccd1 _17050_/Q sky130_fd_sc_hd__dfxtp_1
X_14262_ _15103_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11474_ hold2320/X hold5697/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _13212_/X hold3628/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__mux2_1
X_16001_ _18408_/CLK _16001_/D vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__dfxtp_1
X_10425_ _10998_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__or2_1
X_14193_ hold2170/X _14198_/B _14192_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _13137_/X _13143_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17536_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_104_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10356_ _10548_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13075_ _13074_/X _16902_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__mux2_1
X_17952_ _18071_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
X_10287_ _10557_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__or2_1
X_12026_ hold1108/X hold3353/X _12353_/C vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__mux2_1
X_16903_ _17879_/CLK _16903_/D vssd1 vssd1 vccd1 vccd1 _16903_/Q sky130_fd_sc_hd__dfxtp_1
X_17883_ _17884_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
X_16834_ _18069_/CLK _16834_/D vssd1 vssd1 vccd1 vccd1 _16834_/Q sky130_fd_sc_hd__dfxtp_1
X_16765_ _18025_/CLK _16765_/D vssd1 vssd1 vccd1 vccd1 _16765_/Q sky130_fd_sc_hd__dfxtp_1
X_13977_ hold869/X _13980_/B _13976_/X _13911_/A vssd1 vssd1 vccd1 vccd1 hold870/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15716_ _18426_/CLK _15716_/D vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ hold1140/X _17487_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__mux2_1
X_16696_ _18216_/CLK _16696_/D vssd1 vssd1 vccd1 vccd1 _16696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _18441_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _18445_/CLK _15647_/D vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ hold1263/X _17464_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18366_ _18373_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
X_15578_ _17262_/CLK _15578_/D vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _17318_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 _17317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14529_ _14529_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14529_/X sky130_fd_sc_hd__or2_1
X_18297_ _18330_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08050_ _14218_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _17283_/CLK _17248_/D vssd1 vssd1 vccd1 vccd1 _17248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ _17211_/CLK _17179_/D vssd1 vssd1 vccd1 vccd1 _17179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_321_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17419_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3105 _18112_/Q vssd1 vssd1 vccd1 vccd1 hold3105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3116 _09391_/X vssd1 vssd1 vccd1 vccd1 _16283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3127 _10650_/Y vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08952_ _15414_/A hold320/X vssd1 vssd1 vccd1 vccd1 _16093_/D sky130_fd_sc_hd__and2_1
Xhold3138 _17581_/Q vssd1 vssd1 vccd1 vccd1 hold3138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2404 _14613_/X vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 _12370_/Y vssd1 vssd1 vccd1 vccd1 _17280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _18211_/Q vssd1 vssd1 vccd1 vccd1 hold2415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2426 _08428_/X vssd1 vssd1 vccd1 vccd1 _15844_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07903_ hold2260/X _07924_/B _07902_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07903_/X
+ sky130_fd_sc_hd__o211a_1
X_08883_ _15304_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _16059_/D sky130_fd_sc_hd__and2_1
Xhold2437 _18455_/Q vssd1 vssd1 vccd1 vccd1 hold2437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 _14893_/X vssd1 vssd1 vccd1 vccd1 _18235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _09298_/X vssd1 vssd1 vccd1 vccd1 _16259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _18352_/Q vssd1 vssd1 vccd1 vccd1 hold1714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _18373_/Q vssd1 vssd1 vccd1 vccd1 hold2459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 _18291_/Q vssd1 vssd1 vccd1 vccd1 hold1725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07834_ hold1094/X _07865_/B _07833_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07834_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1736 _15574_/Q vssd1 vssd1 vccd1 vccd1 hold1736/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 _14851_/X vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 _18355_/Q vssd1 vssd1 vccd1 vccd1 hold1758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _15210_/X vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09504_ _09903_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ _07785_/Y hold634/X _15314_/A _09434_/X vssd1 vssd1 vccd1 vccd1 hold635/A
+ sky130_fd_sc_hd__o211a_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09400_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _15541_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_191_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _15519_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__or2_1
XANTENNA_40 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _14972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_62 hold173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _15527_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__or2_1
XANTENNA_73 hold800/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_84 hold5857/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_95 _14545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ _15513_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5030 _17210_/Q vssd1 vssd1 vccd1 vccd1 hold5030/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5041 _09571_/X vssd1 vssd1 vccd1 vccd1 _16347_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10210_ hold4706/X _10568_/B _10209_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5052 _17746_/Q vssd1 vssd1 vccd1 vccd1 hold5052/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11190_ hold5245/X _11121_/A _11189_/X vssd1 vssd1 vccd1 vccd1 _11190_/Y sky130_fd_sc_hd__a21oi_1
Xhold5063 _13756_/X vssd1 vssd1 vccd1 vccd1 _17705_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5074 _17733_/Q vssd1 vssd1 vccd1 vccd1 hold5074/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4340 _11536_/X vssd1 vssd1 vccd1 vccd1 _17002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5085 _10699_/X vssd1 vssd1 vccd1 vccd1 _16723_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10141_ hold3360/X _10619_/B _10140_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _10141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5096 _17062_/Q vssd1 vssd1 vccd1 vccd1 hold5096/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4351 _16606_/Q vssd1 vssd1 vccd1 vccd1 hold4351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4362 _10450_/X vssd1 vssd1 vccd1 vccd1 _16640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4373 _16807_/Q vssd1 vssd1 vccd1 vccd1 hold4373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4384 _13432_/X vssd1 vssd1 vccd1 vccd1 _17597_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4395 _17645_/Q vssd1 vssd1 vccd1 vccd1 hold4395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3650 _11179_/Y vssd1 vssd1 vccd1 vccd1 _16883_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10072_ _10588_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10072_/Y sky130_fd_sc_hd__nor2_1
Xhold3661 _10054_/Y vssd1 vssd1 vccd1 vccd1 _16508_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3672 _13831_/Y vssd1 vssd1 vccd1 vccd1 _17730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3683 _10042_/Y vssd1 vssd1 vccd1 vccd1 _16504_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3694 _10590_/Y vssd1 vssd1 vccd1 vccd1 _10591_/B sky130_fd_sc_hd__dlygate4sd3_1
X_13900_ _15189_/A hold2919/X hold244/X vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__mux2_1
Xhold2960 _14695_/X vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14880_ _15219_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__nand2_1
Xhold2971 _18028_/Q vssd1 vssd1 vccd1 vccd1 hold2971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2982 _15140_/X vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2993 _14514_/X vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13831_ _13864_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16550_ _18118_/CLK _16550_/D vssd1 vssd1 vccd1 vccd1 _16550_/Q sky130_fd_sc_hd__dfxtp_1
X_13762_ hold4567/X _13856_/B _13761_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13762_/X
+ sky130_fd_sc_hd__o211a_1
X_10974_ _11106_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__or2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15517_/A hold1365/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__mux2_1
X_12713_ hold3519/X _12712_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__mux2_1
X_16481_ _18330_/CLK _16481_/D vssd1 vssd1 vccd1 vccd1 _16481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13693_ hold5205/X _13883_/B _13692_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18220_ _18220_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
X_15432_ _15471_/A _15432_/B _15432_/C _15432_/D vssd1 vssd1 vccd1 vccd1 _15432_/X
+ sky130_fd_sc_hd__or4_1
X_12644_ _17391_/Q _12643_/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18151_ _18183_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_15363_ _15481_/A1 _15355_/X _15362_/X _15481_/B1 _18412_/Q vssd1 vssd1 vccd1 vccd1
+ _15363_/X sky130_fd_sc_hd__a32o_1
X_12575_ hold3120/X _12574_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ _17262_/CLK _17102_/D vssd1 vssd1 vccd1 vccd1 _17102_/Q sky130_fd_sc_hd__dfxtp_1
X_14314_ _14529_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14314_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18082_ _18210_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _12204_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__or2_1
X_15294_ _15414_/A _15294_/B vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__and2_1
XFILLER_0_34_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _17882_/CLK _17033_/D vssd1 vssd1 vccd1 vccd1 _17033_/Q sky130_fd_sc_hd__dfxtp_1
X_11457_ _12093_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__or2_1
X_14245_ hold2977/X _14266_/B _14244_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ hold3972/X _10646_/B _10407_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10408_/X
+ sky130_fd_sc_hd__o211a_1
X_14176_ _14246_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14176_/X sky130_fd_sc_hd__or2_1
X_11388_ _11688_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _13183_/A1 _13125_/X _13126_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__o211a_1
X_10339_ hold4061/X _10580_/B _10338_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10339_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _17558_/Q _17092_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__mux2_1
X_17935_ _18033_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_1
X_12009_ _13716_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17866_ _17896_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_1
X_16817_ _18020_/CLK _16817_/D vssd1 vssd1 vccd1 vccd1 _16817_/Q sky130_fd_sc_hd__dfxtp_1
X_17797_ _17829_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16748_ _18241_/CLK _16748_/D vssd1 vssd1 vccd1 vccd1 _16748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16679_ _18205_/CLK _16679_/D vssd1 vssd1 vccd1 vccd1 _16679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _15549_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__or2_1
X_18418_ _18420_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09151_ hold2599/X _09164_/B _09150_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _09151_/X
+ sky130_fd_sc_hd__o211a_1
X_18349_ _18381_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
X_08102_ hold279/X hold606/A hold298/A hold624/A vssd1 vssd1 vccd1 vccd1 hold280/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ hold949/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08033_ _14774_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08033_/Y sky130_fd_sc_hd__nand2_1
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
Xhold800 hold800/A vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__clkbuf_16
Xhold811 hold811/A vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wb_rst_i vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold844 hold844/A vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/A vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 hold866/A vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 la_data_in[23] vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 hold888/A vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 hold926/X vssd1 vssd1 vccd1 vccd1 hold927/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09984_ _09987_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2201 _15788_/Q vssd1 vssd1 vccd1 vccd1 hold2201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2212 _12513_/X vssd1 vssd1 vccd1 vccd1 hold2212/X sky130_fd_sc_hd__dlygate4sd3_1
X_08935_ hold23/X hold456/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08936_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2223 _08032_/X vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2234 _18284_/Q vssd1 vssd1 vccd1 vccd1 hold2234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1500 _14847_/X vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 _15560_/X vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2256 _15563_/Q vssd1 vssd1 vccd1 vccd1 hold2256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 _16223_/Q vssd1 vssd1 vccd1 vccd1 hold1511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2267 _14841_/X vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _14291_/X vssd1 vssd1 vccd1 vccd1 _17945_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08866_ hold291/X hold565/X _08866_/S vssd1 vssd1 vccd1 vccd1 hold566/A sky130_fd_sc_hd__mux2_1
Xhold2278 _14647_/X vssd1 vssd1 vccd1 vccd1 _18116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 _17906_/Q vssd1 vssd1 vccd1 vccd1 hold1533/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1544 _17862_/Q vssd1 vssd1 vccd1 vccd1 hold1544/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2289 _09119_/X vssd1 vssd1 vccd1 vccd1 _16174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 _18222_/Q vssd1 vssd1 vccd1 vccd1 hold1555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 _14803_/X vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ _07817_/A _07817_/B _07817_/C _07817_/D vssd1 vssd1 vccd1 vccd1 _09400_/A
+ sky130_fd_sc_hd__or4_4
X_08797_ hold23/X hold704/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold705/A sky130_fd_sc_hd__mux2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1577 _14901_/X vssd1 vssd1 vccd1 vccd1 _18238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 _15084_/X vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1599 _16205_/Q vssd1 vssd1 vccd1 vccd1 hold1599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _09438_/B _16295_/Q vssd1 vssd1 vccd1 vccd1 _09418_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ hold3974/X _11747_/B _10689_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09349_ _09400_/A _09351_/B _09364_/B vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ hold3819/X _13392_/A _12359_/X vssd1 vssd1 vccd1 vccd1 _12360_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_243_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17708_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ hold5677/X _11789_/B _11310_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _13797_/A _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__or2_1
X_14030_ _15537_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14030_/X sky130_fd_sc_hd__or2_1
X_11242_ hold4619/X _12299_/B _11241_/X _12666_/A vssd1 vssd1 vccd1 vccd1 _11242_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _12331_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11173_/Y sky130_fd_sc_hd__nor2_1
Xhold4170 _13854_/Y vssd1 vssd1 vccd1 vccd1 _13855_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4181 _10510_/X vssd1 vssd1 vccd1 vccd1 _16660_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10124_ hold2683/X hold3132/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__mux2_1
Xhold4192 hold5842/X vssd1 vssd1 vccd1 vccd1 hold5843/A sky130_fd_sc_hd__buf_4
X_15981_ _17300_/CLK _15981_/D vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__dfxtp_1
X_17720_ _17725_/CLK _17720_/D vssd1 vssd1 vccd1 vccd1 _17720_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3480 _10948_/X vssd1 vssd1 vccd1 vccd1 _16806_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3491 _16447_/Q vssd1 vssd1 vccd1 vccd1 hold3491/X sky130_fd_sc_hd__dlygate4sd3_1
X_10055_ _10055_/A _10601_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__and3_1
X_14932_ hold883/X _14964_/B vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2790 _07959_/X vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17651_ _17737_/CLK _17651_/D vssd1 vssd1 vccd1 vccd1 _17651_/Q sky130_fd_sc_hd__dfxtp_1
X_14863_ hold1326/X _14882_/B _14862_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14863_/X
+ sky130_fd_sc_hd__o211a_1
X_16602_ _18224_/CLK _16602_/D vssd1 vssd1 vccd1 vccd1 _16602_/Q sky130_fd_sc_hd__dfxtp_1
X_13814_ _17725_/Q _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13814_/X sky130_fd_sc_hd__and3_1
X_17582_ _17742_/CLK _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
X_14794_ _15187_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16533_ _18219_/CLK _16533_/D vssd1 vssd1 vccd1 vccd1 _16533_/Q sky130_fd_sc_hd__dfxtp_1
X_13745_ hold1426/X _17702_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__mux2_1
X_10957_ hold4091/X _11150_/B _10956_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10957_/X
+ sky130_fd_sc_hd__o211a_1
X_16464_ _18391_/CLK _16464_/D vssd1 vssd1 vccd1 vccd1 _16464_/Q sky130_fd_sc_hd__dfxtp_1
X_13676_ hold2082/X hold3556/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ hold5421/X _11753_/B _10887_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__o211a_1
X_18203_ _18235_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
X_15415_ hold261/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12627_ _12855_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _17385_/D sky130_fd_sc_hd__and2_1
X_16395_ _18380_/CLK _16395_/D vssd1 vssd1 vccd1 vccd1 _16395_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_2__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ _18232_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15346_ _17338_/Q _09362_/C _09362_/D hold528/X vssd1 vssd1 vccd1 vccd1 _15346_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _12924_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _17362_/D sky130_fd_sc_hd__and2_1
XFILLER_0_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11509_ hold4649/X _11798_/B _11508_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11509_/X
+ sky130_fd_sc_hd__o211a_1
X_18065_ _18065_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
X_15277_ hold98/X _09357_/A _15484_/B1 hold222/X _15276_/X vssd1 vssd1 vccd1 vccd1
+ _15282_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12489_ hold8/X _08598_/B _08999_/B _12488_/X _12402_/A vssd1 vssd1 vccd1 vccd1 hold9/A
+ sky130_fd_sc_hd__o311a_1
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold118 hold603/X vssd1 vssd1 vccd1 vccd1 hold604/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__clkbuf_4
X_17016_ _17896_/CLK _17016_/D vssd1 vssd1 vccd1 vccd1 _17016_/Q sky130_fd_sc_hd__dfxtp_1
X_14228_ hold826/X _14230_/B vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ hold2834/X _14148_/B _14158_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout609 _09363_/Y vssd1 vssd1 vccd1 vccd1 _15447_/B1 sky130_fd_sc_hd__buf_8
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _15482_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _15981_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17751_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _18305_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_1
X_08651_ hold65/X hold554/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__mux2_1
X_17849_ _17882_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08582_ hold50/X hold522/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ hold1393/X _09218_/B _09202_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09203_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09134_ _15517_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09065_ _14555_/C hold271/X vssd1 vssd1 vccd1 vccd1 _15508_/B sky130_fd_sc_hd__or2_4
XFILLER_0_13_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08016_ hold2014/X _08029_/B _08015_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _08016_/X
+ sky130_fd_sc_hd__o211a_1
Xhold630 hold630/A vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 la_data_in[31] vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/A vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 hold685/A vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ _10061_/A _10073_/B _09966_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09967_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2020 _15853_/Q vssd1 vssd1 vccd1 vccd1 hold2020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 _09326_/X vssd1 vssd1 vccd1 vccd1 _16273_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2042 _17877_/Q vssd1 vssd1 vccd1 vccd1 hold2042/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ hold251/X hold425/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__mux2_1
Xhold2053 _14436_/X vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _15656_/Q vssd1 vssd1 vccd1 vccd1 hold2064/X sky130_fd_sc_hd__dlygate4sd3_1
X_09898_ hold5683/X _09992_/B _09897_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09898_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _18189_/Q vssd1 vssd1 vccd1 vccd1 hold1330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2075 _15001_/X vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2086 _08212_/X vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 input65/X vssd1 vssd1 vccd1 vccd1 hold1341/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 _14075_/X vssd1 vssd1 vccd1 vccd1 _17842_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 _14339_/X vssd1 vssd1 vccd1 vccd1 _17969_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 _18375_/Q vssd1 vssd1 vccd1 vccd1 hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _15482_/A _08849_/B vssd1 vssd1 vccd1 vccd1 _16043_/D sky130_fd_sc_hd__and2_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _14963_/X vssd1 vssd1 vccd1 vccd1 _18268_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _18285_/Q vssd1 vssd1 vccd1 vccd1 hold1385/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1396 _07996_/X vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ hold5556/X _12338_/B _11859_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11860_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ hold2298/X _16761_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11791_ _11791_/A _11791_/B vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__nor2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13530_ _13734_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10742_ hold2429/X hold5318/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13461_ _13779_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13461_/X sky130_fd_sc_hd__or2_1
X_10673_ hold1016/X hold5294/X _11066_/S vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ hold1290/X _15219_/B _15199_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _15200_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12412_ _12426_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _17299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16180_ _17464_/CLK _16180_/D vssd1 vssd1 vccd1 vccd1 _16180_/Q sky130_fd_sc_hd__dfxtp_1
X_13392_ _13392_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15131_ _15185_/A _15149_/B vssd1 vssd1 vccd1 vccd1 _15131_/X sky130_fd_sc_hd__or2_1
X_12343_ _12343_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _12343_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15062_ _15062_/A _15062_/B vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__and2_1
X_12274_ hold4667/X _12374_/B _12273_/X _12274_/C1 vssd1 vssd1 vccd1 vccd1 _12274_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ hold2505/X _14040_/B _14012_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _14013_/X
+ sky130_fd_sc_hd__o211a_1
X_11225_ _16899_/Q _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ _16876_/Q _11156_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__and3_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ _10491_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15964_ _18425_/CLK _15964_/D vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__dfxtp_1
X_11087_ hold2862/X _16853_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__mux2_1
X_17703_ _17703_/CLK _17703_/D vssd1 vssd1 vccd1 vccd1 _17703_/Q sky130_fd_sc_hd__dfxtp_1
X_10038_ _13214_/A _10098_/A _10037_/X vssd1 vssd1 vccd1 vccd1 _10038_/Y sky130_fd_sc_hd__a21oi_1
X_14915_ hold2559/X _14946_/B _14914_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _14915_/X
+ sky130_fd_sc_hd__o211a_1
X_15895_ _17341_/CLK _15895_/D vssd1 vssd1 vccd1 vccd1 hold533/A sky130_fd_sc_hd__dfxtp_1
X_17634_ _17634_/CLK _17634_/D vssd1 vssd1 vccd1 vccd1 _17634_/Q sky130_fd_sc_hd__dfxtp_1
X_14846_ _15185_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17565_ _17694_/CLK _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ hold766/X _14772_/B _14776_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 hold767/A
+ sky130_fd_sc_hd__o211a_1
X_11989_ hold4710/X _12377_/B _11988_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11989_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16516_ _18236_/CLK _16516_/D vssd1 vssd1 vccd1 vccd1 _16516_/Q sky130_fd_sc_hd__dfxtp_1
X_13728_ _13737_/A _13728_/B vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _17496_/CLK _17496_/D vssd1 vssd1 vccd1 vccd1 _17496_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_165_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18226_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16447_ _18392_/CLK _16447_/D vssd1 vssd1 vccd1 vccd1 _16447_/Q sky130_fd_sc_hd__dfxtp_1
X_13659_ _13788_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16378_ _18355_/CLK _16378_/D vssd1 vssd1 vccd1 vccd1 _16378_/Q sky130_fd_sc_hd__dfxtp_1
X_18117_ _18149_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
X_15329_ _15974_/Q _15485_/A2 _15447_/B1 hold420/X _15328_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/C sky130_fd_sc_hd__a221o_1
Xhold5607 _11059_/X vssd1 vssd1 vccd1 vccd1 _16843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5618 _10675_/X vssd1 vssd1 vccd1 vccd1 _16715_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5629 _16826_/Q vssd1 vssd1 vccd1 vccd1 hold5629/X sky130_fd_sc_hd__dlygate4sd3_1
X_18048_ _18305_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4906 _12106_/X vssd1 vssd1 vccd1 vccd1 _17192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4917 _17209_/Q vssd1 vssd1 vccd1 vccd1 hold4917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4928 _11623_/X vssd1 vssd1 vccd1 vccd1 _17031_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4939 _16993_/Q vssd1 vssd1 vccd1 vccd1 hold4939/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout406 _14334_/B vssd1 vssd1 vccd1 vccd1 _14338_/B sky130_fd_sc_hd__clkbuf_8
X_09821_ hold2372/X _16431_/Q _10028_/C vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__mux2_1
Xfanout417 hold586/X vssd1 vssd1 vccd1 vccd1 hold587/A sky130_fd_sc_hd__buf_1
Xfanout428 hold243/X vssd1 vssd1 vccd1 vccd1 _13942_/S sky130_fd_sc_hd__buf_4
Xfanout439 _12308_/C vssd1 vssd1 vccd1 vccd1 _13796_/S sky130_fd_sc_hd__buf_6
X_09752_ hold2196/X _16408_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08703_ hold17/X hold221/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__mux2_1
X_09683_ hold1348/X hold3484/X _10628_/C vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _15414_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _15939_/D sky130_fd_sc_hd__and2_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08970_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _15906_/D sky130_fd_sc_hd__and2_1
X_08496_ _14728_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ hold2945/X _09119_/A2 _09116_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09117_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ hold251/X hold375/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold471 hold471/A vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 hold482/A vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _11106_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout940 _14866_/A vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__clkbuf_8
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ hold2851/X hold3073/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__mux2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _15034_/X vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14986_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14700_/X sky130_fd_sc_hd__or2_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 _17974_/Q vssd1 vssd1 vccd1 vccd1 hold1171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _14931_/X vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ hold1677/X _17128_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__mux2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _17897_/CLK _15680_/D vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _15706_/Q vssd1 vssd1 vccd1 vccd1 hold1193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ hold1185/X _17475_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__mux2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ hold1732/X _14666_/B _14630_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _14631_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ hold2766/X hold3835/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17513_/CLK _17350_/D vssd1 vssd1 vccd1 vccd1 _17350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _15492_/A _14573_/B hold1794/X vssd1 vssd1 vccd1 vccd1 _14562_/X sky130_fd_sc_hd__a21o_1
X_11774_ _11774_/A _12338_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and3_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _17503_/CLK hold682/X vssd1 vssd1 vccd1 vccd1 _16301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13513_ hold3212/X _13808_/B _13512_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13513_/X
+ sky130_fd_sc_hd__o211a_1
X_17281_ _17281_/CLK _17281_/D vssd1 vssd1 vccd1 vccd1 _17281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _11667_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__or2_1
X_14493_ hold770/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14493_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16232_ _17435_/CLK _16232_/D vssd1 vssd1 vccd1 vccd1 hold997/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ hold4465/X _13832_/B _13443_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13444_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _11136_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16163_ _18013_/CLK _16163_/D vssd1 vssd1 vccd1 vccd1 _16163_/Q sky130_fd_sc_hd__dfxtp_1
X_10587_ _16526_/Q _09951_/A _10586_/X vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13375_ hold5164/X _13883_/B _13374_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13375_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ hold2100/X _15113_/B _15113_/Y _15058_/A vssd1 vssd1 vccd1 vccd1 _15114_/X
+ sky130_fd_sc_hd__o211a_1
X_12326_ _17266_/Q _13871_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__and3_1
X_16094_ _17302_/CLK _16094_/D vssd1 vssd1 vccd1 vccd1 hold495/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ _15099_/A hold2643/X hold302/X vssd1 vssd1 vccd1 vccd1 _15046_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ hold2291/X _17243_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ hold5447/X _11694_/A _11207_/X vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__a21oi_1
X_12188_ hold1834/X hold4729/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__mux2_1
X_11139_ _11637_/A _11139_/B vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__or2_1
X_16996_ _17844_/CLK _16996_/D vssd1 vssd1 vccd1 vccd1 _16996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ _17329_/CLK _15947_/D vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15878_ _17749_/CLK _15878_/D vssd1 vssd1 vccd1 vccd1 _15878_/Q sky130_fd_sc_hd__dfxtp_1
X_17617_ _17649_/CLK _17617_/D vssd1 vssd1 vccd1 vccd1 _17617_/Q sky130_fd_sc_hd__dfxtp_1
X_14829_ hold1152/X _14828_/B _14828_/Y _15072_/A vssd1 vssd1 vccd1 vccd1 _14829_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08350_ _14854_/A hold2383/X hold122/X vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__mux2_1
X_17548_ _18185_/CLK _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08281_ hold2024/X _08268_/B _08280_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _08281_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _17480_/CLK _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5404 _11470_/X vssd1 vssd1 vccd1 vccd1 _16980_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5415 _16465_/Q vssd1 vssd1 vccd1 vccd1 hold5415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5426 _09541_/X vssd1 vssd1 vccd1 vccd1 _16337_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5437 _16428_/Q vssd1 vssd1 vccd1 vccd1 hold5437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4703 _11608_/X vssd1 vssd1 vccd1 vccd1 _17026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5448 _11208_/Y vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4714 _16691_/Q vssd1 vssd1 vccd1 vccd1 hold4714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5459 _09817_/X vssd1 vssd1 vccd1 vccd1 _16429_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4725 _17007_/Q vssd1 vssd1 vccd1 vccd1 hold4725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4736 _10276_/X vssd1 vssd1 vccd1 vccd1 _16582_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4747 _17744_/Q vssd1 vssd1 vccd1 vccd1 hold4747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4758 _10894_/X vssd1 vssd1 vccd1 vccd1 _16788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4769 _17129_/Q vssd1 vssd1 vccd1 vccd1 hold4769/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout203 _11792_/B vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__buf_4
Xfanout214 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10780_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout225 _10465_/A2 vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__buf_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 _09952_/A2 vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__buf_4
Xfanout247 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__clkbuf_4
X_09804_ _09903_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__or2_1
Xfanout258 fanout299/X vssd1 vssd1 vccd1 vccd1 _13674_/A sky130_fd_sc_hd__buf_2
Xfanout269 fanout299/X vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__buf_2
X_07996_ hold1395/X _08029_/B _07995_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07996_/X
+ sky130_fd_sc_hd__o211a_1
X_09735_ _10560_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ _09975_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__or2_1
X_08617_ hold443/X hold643/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08618_/B sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09987_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__or2_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ hold126/X hold373/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08479_ hold808/X _08486_/B _08478_/X _08381_/A vssd1 vssd1 vccd1 vccd1 hold809/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ hold4180/X _10589_/B _10509_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10510_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11490_ _12093_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ hold4147/X _10631_/B _10440_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ _13153_/X _13159_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17538_/D sky130_fd_sc_hd__o21a_1
X_10372_ hold3554/X _10558_/A2 _10371_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10372_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _13716_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__or2_1
X_13091_ _13090_/X _16904_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
Xhold5960 _18048_/Q vssd1 vssd1 vccd1 vccd1 hold5960/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5971 _18036_/Q vssd1 vssd1 vccd1 vccd1 hold5971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5982 _18369_/Q vssd1 vssd1 vccd1 vccd1 hold5982/X sky130_fd_sc_hd__dlygate4sd3_1
X_12042_ _12234_/A _12042_/B vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__or2_1
Xhold5993 _18415_/Q vssd1 vssd1 vccd1 vccd1 hold5993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 input29/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__buf_1
X_16850_ _18053_/CLK _16850_/D vssd1 vssd1 vccd1 vccd1 _16850_/Q sky130_fd_sc_hd__dfxtp_1
X_15801_ _17669_/CLK _15801_/D vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout770 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _12256_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout781 _14388_/A vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__buf_4
X_16781_ _17984_/CLK _16781_/D vssd1 vssd1 vccd1 vccd1 _16781_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout792 _15056_/A vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__buf_4
X_13993_ hold2193/X _13980_/B _13992_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _13993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _17703_/CLK _15732_/D vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfxtp_1
X_12944_ hold3587/X _12943_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__mux2_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18451_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
X_15663_ _17216_/CLK _15663_/D vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ hold3109/X _12874_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__mux2_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _18454_/CLK _17402_/D vssd1 vssd1 vccd1 vccd1 _17402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _15169_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18382_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
X_11826_ _12018_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__or2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _17274_/CLK _15594_/D vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _18410_/CLK hold185/X vssd1 vssd1 vccd1 vccd1 _17333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _15225_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14545_/X sky130_fd_sc_hd__or2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ hold5227/X _11667_/A _11756_/X vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _17844_/CLK _17264_/D vssd1 vssd1 vccd1 vccd1 _17264_/Q sky130_fd_sc_hd__dfxtp_1
X_10708_ hold4591/X _11192_/B _10707_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14476_ hold1748/X _14481_/B _14475_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14476_/X
+ sky130_fd_sc_hd__o211a_1
X_11688_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11688_/X sky130_fd_sc_hd__or2_1
X_16215_ _17447_/CLK _16215_/D vssd1 vssd1 vccd1 vccd1 _16215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13427_ hold2513/X hold4828/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__mux2_1
X_10639_ _10651_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__nor2_1
X_17195_ _17227_/CLK _17195_/D vssd1 vssd1 vccd1 vccd1 _17195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ _17341_/CLK _16146_/D vssd1 vssd1 vccd1 vccd1 hold642/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13358_ hold1225/X hold3846/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12309_ hold3141/X _12210_/A _12308_/X vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16077_ _18405_/CLK _16077_/D vssd1 vssd1 vccd1 vccd1 hold425/A sky130_fd_sc_hd__dfxtp_1
X_13289_ _13289_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__and2_1
Xhold3309 _17463_/Q vssd1 vssd1 vccd1 vccd1 hold3309/X sky130_fd_sc_hd__dlygate4sd3_1
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__and2_1
Xhold2608 _14021_/X vssd1 vssd1 vccd1 vccd1 _17816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2619 _14969_/X vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07850_ hold2220/X _07869_/B _07849_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07850_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1907 _16186_/Q vssd1 vssd1 vccd1 vccd1 hold1907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 _09167_/X vssd1 vssd1 vccd1 vccd1 _16196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1929 _15816_/Q vssd1 vssd1 vccd1 vccd1 hold1929/X sky130_fd_sc_hd__dlygate4sd3_1
X_07781_ hold335/X vssd1 vssd1 vccd1 vccd1 _07781_/Y sky130_fd_sc_hd__inv_2
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _17891_/CLK _16979_/D vssd1 vssd1 vccd1 vccd1 _16979_/Q sky130_fd_sc_hd__dfxtp_1
X_09520_ hold5598/X _09998_/B _09519_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09520_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_180_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ _09456_/C _09456_/D _09450_/Y vssd1 vssd1 vccd1 vccd1 _16310_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ hold1640/X _08440_/A2 _08401_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _08402_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ hold717/X _09392_/B _09362_/D hold670/X _09381_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _15557_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _15543_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08195_ _15529_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5201 _17674_/Q vssd1 vssd1 vccd1 vccd1 hold5201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5212 _13786_/X vssd1 vssd1 vccd1 vccd1 _17715_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5223 _10015_/Y vssd1 vssd1 vccd1 vccd1 _16495_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5234 _11754_/Y vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4500 _17694_/Q vssd1 vssd1 vccd1 vccd1 hold4500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5245 _16727_/Q vssd1 vssd1 vccd1 vccd1 hold5245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4511 _10411_/X vssd1 vssd1 vccd1 vccd1 _16627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5256 _11176_/Y vssd1 vssd1 vccd1 vccd1 _16882_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4522 _16373_/Q vssd1 vssd1 vccd1 vccd1 hold4522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5267 _11214_/Y vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5278 _17110_/Q vssd1 vssd1 vccd1 vccd1 hold5278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4533 _11647_/X vssd1 vssd1 vccd1 vccd1 _17039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4544 _17588_/Q vssd1 vssd1 vccd1 vccd1 hold4544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5289 _16922_/Q vssd1 vssd1 vccd1 vccd1 hold5289/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3810 _12304_/Y vssd1 vssd1 vccd1 vccd1 _17258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4555 _16997_/Q vssd1 vssd1 vccd1 vccd1 hold4555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4566 _10387_/X vssd1 vssd1 vccd1 vccd1 _16619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3821 _12361_/Y vssd1 vssd1 vccd1 vccd1 _17277_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3832 _09523_/X vssd1 vssd1 vccd1 vccd1 _16331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4577 _16009_/Q vssd1 vssd1 vccd1 vccd1 _15395_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3843 _11800_/Y vssd1 vssd1 vccd1 vccd1 _17090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4588 _10777_/X vssd1 vssd1 vccd1 vccd1 _16749_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3854 _10585_/Y vssd1 vssd1 vccd1 vccd1 _16685_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4599 _17180_/Q vssd1 vssd1 vccd1 vccd1 hold4599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3865 _17562_/Q vssd1 vssd1 vccd1 vccd1 hold3865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3876 _10588_/Y vssd1 vssd1 vccd1 vccd1 _16686_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_268_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17170_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3887 _10918_/X vssd1 vssd1 vccd1 vccd1 _16796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3898 _12357_/Y vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07979_ hold1861/X _07978_/B _07978_/Y _08163_/A vssd1 vssd1 vccd1 vccd1 _07979_/X
+ sky130_fd_sc_hd__o211a_1
X_09718_ hold5437/X _10013_/B _09717_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__o211a_1
X_10990_ hold4721/X _11192_/B _10989_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09649_ hold3283/X _09952_/A2 _09648_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09649_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _15502_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _17396_/D sky130_fd_sc_hd__and2_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ hold4967/X _11792_/B _11610_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11611_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _15506_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _17373_/D sky130_fd_sc_hd__and2_1
XFILLER_0_132_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14330_ _14330_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14330_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ hold4813/X _11732_/B _11541_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ hold1704/X _14266_/B _14260_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14261_/X
+ sky130_fd_sc_hd__o211a_1
X_11473_ hold5731/X _11789_/B _11472_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16000_ _18407_/CLK _16000_/D vssd1 vssd1 vccd1 vccd1 hold632/A sky130_fd_sc_hd__dfxtp_1
X_13212_ hold5245/X _13211_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_2
X_10424_ hold2995/X _16632_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__mux2_1
X_14192_ _15537_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14192_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13143_ _13183_/A1 _13141_/X _13142_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13143_/X
+ sky130_fd_sc_hd__o211a_1
X_10355_ hold2807/X _16609_/Q _10643_/C vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__mux2_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5790 hold5790/A vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_12
X_13074_ _17560_/Q _17094_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _18241_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
X_10286_ hold2938/X hold3533/X _10562_/S vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__mux2_1
X_12025_ hold4965/X _12311_/B _12024_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _12025_/X
+ sky130_fd_sc_hd__o211a_1
X_16902_ _18428_/CLK _16902_/D vssd1 vssd1 vccd1 vccd1 _16902_/Q sky130_fd_sc_hd__dfxtp_1
X_17882_ _17882_/CLK hold970/X vssd1 vssd1 vccd1 vccd1 hold969/A sky130_fd_sc_hd__dfxtp_1
X_16833_ _18070_/CLK _16833_/D vssd1 vssd1 vccd1 vccd1 _16833_/Q sky130_fd_sc_hd__dfxtp_1
X_16764_ _18060_/CLK _16764_/D vssd1 vssd1 vccd1 vccd1 _16764_/Q sky130_fd_sc_hd__dfxtp_1
X_13976_ hold735/X _13992_/B vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15715_ _17281_/CLK _15715_/D vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12927_ _12927_/A _12927_/B vssd1 vssd1 vccd1 vccd1 _17485_/D sky130_fd_sc_hd__and2_1
X_16695_ _18221_/CLK _16695_/D vssd1 vssd1 vccd1 vccd1 _16695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ _17128_/CLK _15646_/D vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_18434_ _18441_/CLK hold996/X vssd1 vssd1 vccd1 vccd1 hold995/A sky130_fd_sc_hd__dfxtp_1
X_12858_ _12924_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _17462_/D sky130_fd_sc_hd__and2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18365_ _18373_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
X_11809_ hold4379/X _12308_/B _11808_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _11809_/X
+ sky130_fd_sc_hd__o211a_1
X_15577_ _17743_/CLK _15577_/D vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12789_ _12789_/A _12789_/B vssd1 vssd1 vccd1 vccd1 _17439_/D sky130_fd_sc_hd__and2_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17523_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _17316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ hold2754/X _14554_/A2 _14527_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14528_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18296_ _18392_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _17279_/CLK _17247_/D vssd1 vssd1 vccd1 vccd1 _17247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14459_ _15193_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ _17274_/CLK _17178_/D vssd1 vssd1 vccd1 vccd1 _17178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _17524_/CLK _16129_/D vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3106 _14639_/X vssd1 vssd1 vccd1 vccd1 _18112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3117 hold5868/X vssd1 vssd1 vccd1 vccd1 hold5869/A sky130_fd_sc_hd__buf_4
X_08951_ hold126/X _16093_/Q _08993_/S vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__mux2_1
Xhold3128 _10651_/Y vssd1 vssd1 vccd1 vccd1 _16707_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 _13863_/Y vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2405 _18099_/Q vssd1 vssd1 vccd1 vccd1 hold2405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2416 _14845_/X vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07902_ _15525_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07902_/X sky130_fd_sc_hd__or2_1
Xhold2427 _17967_/Q vssd1 vssd1 vccd1 vccd1 hold2427/X sky130_fd_sc_hd__dlygate4sd3_1
X_08882_ hold26/X hold576/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__mux2_1
Xhold2438 _15554_/X vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _15645_/Q vssd1 vssd1 vccd1 vccd1 hold2449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 _17931_/Q vssd1 vssd1 vccd1 vccd1 hold1704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1715 _15138_/X vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1726 _15011_/X vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ hold756/X _07881_/B vssd1 vssd1 vccd1 vccd1 _07833_/X sky130_fd_sc_hd__or2_1
Xhold1737 _07858_/X vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1748 _18035_/Q vssd1 vssd1 vccd1 vccd1 hold1748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1759 _15144_/X vssd1 vssd1 vccd1 vccd1 _18355_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09503_ hold1576/X _16325_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09434_ hold616/X _16303_/Q vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09365_ _09386_/A _09365_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09369_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_191_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08316_ hold1041/X _08323_/B _08315_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08316_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09296_ hold1172/X _09338_/A2 _09295_/X _12927_/A vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_30 _09494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_41 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _14972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_63 hold335/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ hold2534/X _08268_/B _08246_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08247_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_74 hold800/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_85 hold5857/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _14545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08178_ hold922/X _08209_/B _08177_/X _08371_/A vssd1 vssd1 vccd1 vccd1 hold923/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5020 _12160_/X vssd1 vssd1 vccd1 vccd1 _17210_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5031 _12064_/X vssd1 vssd1 vccd1 vccd1 _17178_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5042 _17133_/Q vssd1 vssd1 vccd1 vccd1 hold5042/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5053 _13783_/X vssd1 vssd1 vccd1 vccd1 _17714_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5064 _16961_/Q vssd1 vssd1 vccd1 vccd1 hold5064/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5075 _13744_/X vssd1 vssd1 vccd1 vccd1 _17701_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4330 _09772_/X vssd1 vssd1 vccd1 vccd1 _16414_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10140_ _10524_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__or2_1
Xhold4341 _16774_/Q vssd1 vssd1 vccd1 vccd1 hold4341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5086 _17607_/Q vssd1 vssd1 vccd1 vccd1 hold5086/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5097 _11620_/X vssd1 vssd1 vccd1 vccd1 _17030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4352 _10252_/X vssd1 vssd1 vccd1 vccd1 _16574_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4363 _16865_/Q vssd1 vssd1 vccd1 vccd1 hold4363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4374 _10855_/X vssd1 vssd1 vccd1 vccd1 _16775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3640 _10626_/Y vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4385 _17665_/Q vssd1 vssd1 vccd1 vccd1 hold4385/X sky130_fd_sc_hd__dlygate4sd3_1
X_10071_ _13302_/A _09975_/A _10070_/X vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__a21oi_1
Xhold4396 _13480_/X vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3651 _17569_/Q vssd1 vssd1 vccd1 vccd1 hold3651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3662 _16521_/Q vssd1 vssd1 vccd1 vccd1 hold3662/X sky130_fd_sc_hd__clkbuf_2
Xhold3673 _16522_/Q vssd1 vssd1 vccd1 vccd1 hold3673/X sky130_fd_sc_hd__clkbuf_2
Xhold3684 _16543_/Q vssd1 vssd1 vccd1 vccd1 hold3684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3695 _10591_/Y vssd1 vssd1 vccd1 vccd1 _16687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2950 _14408_/X vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2961 _15830_/Q vssd1 vssd1 vccd1 vccd1 hold2961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2972 _14462_/X vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2983 _18249_/Q vssd1 vssd1 vccd1 vccd1 hold2983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2994 _15693_/Q vssd1 vssd1 vccd1 vccd1 hold2994/X sky130_fd_sc_hd__dlygate4sd3_1
X_13830_ _17570_/Q _13734_/A _13829_/X vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13776_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__or2_1
X_10973_ _18018_/Q hold5719/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__mux2_1
X_15500_ _15502_/A _15500_/B vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__and2_1
X_12712_ hold1107/X hold3497/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16480_ _18235_/CLK _16480_/D vssd1 vssd1 vccd1 vccd1 _16480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13788_/A _13692_/B vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15431_ hold326/X _15451_/A2 _09386_/D hold524/X _15426_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ hold1846/X _17392_/Q _12679_/S vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ _18214_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_1__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_6_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15362_ _15471_/A _15362_/B _15362_/C _15362_/D vssd1 vssd1 vccd1 vccd1 _15362_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_38_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12574_ hold1781/X hold3076/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17101_ _17718_/CLK _17101_/D vssd1 vssd1 vccd1 vccd1 _17101_/Q sky130_fd_sc_hd__dfxtp_1
X_14313_ hold1443/X _14333_/A2 _14312_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _14313_/X
+ sky130_fd_sc_hd__o211a_1
X_18081_ _18392_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
X_11525_ hold2330/X hold4700/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15293_ _15490_/A1 _15285_/X _15292_/X _15490_/B1 hold5841/A vssd1 vssd1 vccd1 vccd1
+ _15293_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17032_ _17880_/CLK _17032_/D vssd1 vssd1 vccd1 vccd1 _17032_/Q sky130_fd_sc_hd__dfxtp_1
X_14244_ _15193_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ hold1799/X hold4441/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _10521_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ hold2909/X _14198_/B _14174_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__o211a_1
X_11387_ hold760/X _16953_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _13126_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__or2_1
X_10338_ _10485_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13055_/C _13057_/B _17521_/Q vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__and3b_4
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _18391_/CLK hold933/X vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10269_ _11097_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12008_ hold2626/X _17160_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__mux2_1
X_17865_ _17865_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16816_ _18052_/CLK _16816_/D vssd1 vssd1 vccd1 vccd1 _16816_/Q sky130_fd_sc_hd__dfxtp_1
X_17796_ _17862_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13959_ hold904/X _13980_/B _13958_/X _15506_/A vssd1 vssd1 vccd1 vccd1 hold905/A
+ sky130_fd_sc_hd__o211a_1
X_16747_ _18305_/CLK _16747_/D vssd1 vssd1 vccd1 vccd1 _16747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ _18236_/CLK _16678_/D vssd1 vssd1 vccd1 vccd1 _16678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18417_ _18417_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15629_ _17257_/CLK _15629_/D vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09150_ _15533_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__or2_1
X_18348_ _18380_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08101_ hold2207/X _08088_/B _08100_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _18424_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ hold2826/X _09119_/A2 _09080_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08032_ hold2222/X _08033_/B _08031_/Y _13933_/A vssd1 vssd1 vccd1 vccd1 _08032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 input50/A vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_6
XFILLER_0_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold801 hold801/A vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 la_data_in[30] vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold834 hold834/A vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 hold845/A vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 hold856/A vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 hold878/A vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ hold2957/X hold5664/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__mux2_1
Xhold889 hold889/A vssd1 vssd1 vccd1 vccd1 input48/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2202 _08310_/X vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _08934_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _08965_/S sky130_fd_sc_hd__or2_2
Xhold2213 _12679_/S vssd1 vssd1 vccd1 vccd1 _12589_/S sky130_fd_sc_hd__clkbuf_4
Xhold2224 _17392_/Q vssd1 vssd1 vccd1 vccd1 hold2224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 _14997_/X vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1501 _15765_/Q vssd1 vssd1 vccd1 vccd1 hold1501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 _18042_/Q vssd1 vssd1 vccd1 vccd1 hold2246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _09223_/X vssd1 vssd1 vccd1 vccd1 _16223_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ _15050_/A hold111/X vssd1 vssd1 vccd1 vccd1 _16051_/D sky130_fd_sc_hd__and2_1
Xhold2257 _07836_/X vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _18324_/Q vssd1 vssd1 vccd1 vccd1 hold1523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 _18152_/Q vssd1 vssd1 vccd1 vccd1 hold2268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2279 _15873_/Q vssd1 vssd1 vccd1 vccd1 hold2279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _14207_/X vssd1 vssd1 vccd1 vccd1 _17906_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1545 _14117_/X vssd1 vssd1 vccd1 vccd1 _17862_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1556 _14867_/X vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ _15515_/A _14972_/A hold892/A _15183_/A vssd1 vssd1 vccd1 vccd1 _07817_/D
+ sky130_fd_sc_hd__or4_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 _18330_/Q vssd1 vssd1 vccd1 vccd1 hold1567/X sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ _08868_/B _08934_/A _13046_/D vssd1 vssd1 vccd1 vccd1 _08801_/S sky130_fd_sc_hd__or3_2
Xhold1578 hold6019/X vssd1 vssd1 vccd1 vccd1 _09463_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1589 _18349_/Q vssd1 vssd1 vccd1 vccd1 hold1589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09417_ _07804_/A _09456_/A _15304_/A _09416_/X vssd1 vssd1 vccd1 vccd1 _09417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ hold86/X _15541_/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09279_ hold800/X hold2678/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11310_ _11694_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11310_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ hold2254/X hold4267/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ _11616_/A _11241_/B vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_283_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17855_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ hold3129/X _11076_/A _11171_/X vssd1 vssd1 vccd1 vccd1 _11172_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_212_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17798_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4160 _10987_/X vssd1 vssd1 vccd1 vccd1 _16819_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10123_ hold5011/X _10073_/B _10122_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10123_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4171 _13855_/Y vssd1 vssd1 vccd1 vccd1 _17738_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4182 _16642_/Q vssd1 vssd1 vccd1 vccd1 hold4182/X sky130_fd_sc_hd__dlygate4sd3_1
X_15980_ _18414_/CLK _15980_/D vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__dfxtp_1
Xhold4193 _15323_/X vssd1 vssd1 vccd1 vccd1 _15324_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3470 _17204_/Q vssd1 vssd1 vccd1 vccd1 hold3470/X sky130_fd_sc_hd__dlygate4sd3_1
X_14931_ hold1181/X _14946_/B _14930_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _14931_/X
+ sky130_fd_sc_hd__o211a_1
X_10054_ _10588_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10054_/Y sky130_fd_sc_hd__nor2_1
Xhold3481 _17353_/Q vssd1 vssd1 vccd1 vccd1 hold3481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3492 _09775_/X vssd1 vssd1 vccd1 vccd1 _16415_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2780 _13048_/X vssd1 vssd1 vccd1 vccd1 _17525_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14862_ hold883/X _14894_/B vssd1 vssd1 vccd1 vccd1 _14862_/X sky130_fd_sc_hd__or2_1
Xhold2791 _15733_/Q vssd1 vssd1 vccd1 vccd1 hold2791/X sky130_fd_sc_hd__dlygate4sd3_1
X_17650_ _17747_/CLK _17650_/D vssd1 vssd1 vccd1 vccd1 _17650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16601_ _18223_/CLK _16601_/D vssd1 vssd1 vccd1 vccd1 _16601_/Q sky130_fd_sc_hd__dfxtp_1
X_13813_ _13822_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__nor2_1
X_17581_ _17741_/CLK _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14793_ hold1489/X _14822_/B _14792_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14793_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16532_ _18218_/CLK _16532_/D vssd1 vssd1 vccd1 vccd1 _16532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ hold5074/X _13856_/B _13743_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _11061_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16463_ _18381_/CLK _16463_/D vssd1 vssd1 vccd1 vccd1 _16463_/Q sky130_fd_sc_hd__dfxtp_1
X_13675_ hold3416/X _13823_/B _13674_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13675_/X
+ sky130_fd_sc_hd__o211a_1
X_10887_ _11658_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__or2_1
X_15414_ _15414_/A _15414_/B vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18202_ _18204_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
X_12626_ hold3078/X _12625_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__mux2_1
X_16394_ _18371_/CLK _16394_/D vssd1 vssd1 vccd1 vccd1 _16394_/Q sky130_fd_sc_hd__dfxtp_1
X_18133_ _18183_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15345_ hold720/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15345_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ hold3244/X _12556_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11508_ _11697_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11508_/X sky130_fd_sc_hd__or2_1
X_18064_ _18064_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_15276_ _17331_/Q _15486_/B1 _15485_/B1 hold199/X vssd1 vssd1 vccd1 vccd1 _15276_/X
+ sky130_fd_sc_hd__a22o_1
X_12488_ _17337_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold584/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17895_/CLK _17015_/D vssd1 vssd1 vccd1 vccd1 _17015_/Q sky130_fd_sc_hd__dfxtp_1
Xhold119 hold605/X vssd1 vssd1 vccd1 vccd1 hold606/A sky130_fd_sc_hd__buf_4
X_14227_ hold1461/X _14216_/Y _14226_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14227_/X
+ sky130_fd_sc_hd__o211a_1
X_11439_ _11631_/A _11439_/B vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14158_ _15557_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14158_/X sky130_fd_sc_hd__or2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13108_/X hold3673/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__mux2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ hold1998/X _14094_/B _14088_/Y _15504_/A vssd1 vssd1 vccd1 vccd1 _14089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _18042_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_1
X_08650_ _12402_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _15947_/D sky130_fd_sc_hd__and2_1
X_17848_ _17877_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_1
X_08581_ _12428_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _15914_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_87_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17318_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _17779_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _15531_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09133_ hold1619/X _09177_/A2 _09132_/X _12924_/A vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09064_ _18461_/Q hold270/X vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08015_ _15529_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_170_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 hold620/A vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold631 hold631/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 hold642/A vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 hold653/A vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 hold664/A vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 hold686/A vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 hold697/A vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _10098_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__or2_1
Xhold2010 _15603_/Q vssd1 vssd1 vccd1 vccd1 hold2010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _08446_/X vssd1 vssd1 vccd1 vccd1 _15853_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08917_ _12428_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _16076_/D sky130_fd_sc_hd__and2_1
Xhold2032 _15741_/Q vssd1 vssd1 vccd1 vccd1 hold2032/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 _14147_/X vssd1 vssd1 vccd1 vccd1 _17877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2054 _17858_/Q vssd1 vssd1 vccd1 vccd1 hold2054/X sky130_fd_sc_hd__dlygate4sd3_1
X_09897_ _11067_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__or2_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2065 _08030_/X vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1320 _17897_/Q vssd1 vssd1 vccd1 vccd1 hold1320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _14799_/X vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2076 _15597_/Q vssd1 vssd1 vccd1 vccd1 hold2076/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _15195_/X vssd1 vssd1 vccd1 vccd1 hold1342/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ hold140/X hold507/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08849_/B sky130_fd_sc_hd__mux2_1
Xhold2087 _16242_/Q vssd1 vssd1 vccd1 vccd1 hold2087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2098 _18365_/Q vssd1 vssd1 vccd1 vccd1 hold2098/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 _17854_/Q vssd1 vssd1 vccd1 vccd1 hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 _15186_/X vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _15628_/Q vssd1 vssd1 vccd1 vccd1 hold1375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 _14999_/X vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ hold251/X _16010_/Q _08787_/S vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__mux2_1
Xhold1397 _15865_/Q vssd1 vssd1 vccd1 vccd1 hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ hold5657/X _11213_/B _10809_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10810_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ hold5321/X _11694_/A _11789_/X vssd1 vssd1 vccd1 vccd1 _11790_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ hold4211/X _11765_/B _10740_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _10741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ hold2425/X _17607_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10672_ hold5490/X _11150_/B _10671_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ hold179/X hold596/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ hold2279/X hold3945/X _13871_/C vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15130_ hold2390/X _15161_/B _15129_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _15130_/X
+ sky130_fd_sc_hd__o211a_1
X_12342_ hold3877/X _12246_/A _12341_/X vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _15169_/A hold1893/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15062_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _12282_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__or2_1
X_14012_ _15519_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__or2_1
X_11224_ _12343_/A _11224_/B vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11155_ _11155_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__nor2_1
X_10106_ hold2893/X _16526_/Q _10628_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__mux2_1
X_15963_ _17318_/CLK _15963_/D vssd1 vssd1 vccd1 vccd1 hold672/A sky130_fd_sc_hd__dfxtp_1
X_11086_ hold4645/X _11192_/B _11085_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _11086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17702_ _17734_/CLK _17702_/D vssd1 vssd1 vccd1 vccd1 _17702_/Q sky130_fd_sc_hd__dfxtp_1
X_14914_ _15129_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14914_/X sky130_fd_sc_hd__or2_1
X_10037_ _16503_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__and3_1
X_15894_ _17340_/CLK _15894_/D vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17633_ _17697_/CLK _17633_/D vssd1 vssd1 vccd1 vccd1 _17633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14845_ hold2415/X _14880_/B _14844_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14776_ hold730/X _14786_/B vssd1 vssd1 vccd1 vccd1 _14776_/X sky130_fd_sc_hd__or2_1
X_17564_ _17724_/CLK _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_1
X_11988_ _12282_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16515_ _18388_/CLK _16515_/D vssd1 vssd1 vccd1 vccd1 _16515_/Q sky130_fd_sc_hd__dfxtp_1
X_13727_ hold922/X hold4325/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13728_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_156_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10939_ hold5661/X _11765_/B _10938_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _16803_/D
+ sky130_fd_sc_hd__o211a_1
X_17495_ _17496_/CLK _17495_/D vssd1 vssd1 vccd1 vccd1 _17495_/Q sky130_fd_sc_hd__dfxtp_1
X_13658_ hold1335/X hold3560/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16446_ _18391_/CLK _16446_/D vssd1 vssd1 vccd1 vccd1 _16446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ _12909_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _17379_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16377_ _18358_/CLK _16377_/D vssd1 vssd1 vccd1 vccd1 _16377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ hold1027/X _17650_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ _18265_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
X_15328_ hold511/X _15484_/A2 _15451_/A2 hold589/X vssd1 vssd1 vccd1 vccd1 _15328_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18386_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5608 _16845_/Q vssd1 vssd1 vccd1 vccd1 hold5608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5619 _16510_/Q vssd1 vssd1 vccd1 vccd1 hold5619/X sky130_fd_sc_hd__dlygate4sd3_1
X_15259_ hold701/X _15485_/A2 _15447_/B1 _16030_/Q _15258_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18047_ _18047_/CLK hold896/X vssd1 vssd1 vccd1 vccd1 hold895/A sky130_fd_sc_hd__dfxtp_1
Xhold4907 _17594_/Q vssd1 vssd1 vccd1 vccd1 hold4907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4918 _12061_/X vssd1 vssd1 vccd1 vccd1 _17177_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4929 _17091_/Q vssd1 vssd1 vccd1 vccd1 hold4929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ hold3711/X _10028_/B _09819_/X _15364_/A vssd1 vssd1 vccd1 vccd1 _09820_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout407 _14286_/Y vssd1 vssd1 vccd1 vccd1 _14333_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout418 _14072_/B vssd1 vssd1 vccd1 vccd1 _14106_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout429 _13056_/X vssd1 vssd1 vccd1 vccd1 _13251_/S sky130_fd_sc_hd__buf_8
X_09751_ hold4607/X _10049_/B _09750_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08702_ _15314_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _15972_/D sky130_fd_sc_hd__and2_1
X_09682_ hold3398/X _10067_/B _09681_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _09682_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08633_ hold184/X hold460/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ hold214/X hold518/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08565_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08495_ hold1866/X _08486_/B _08494_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _08495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ _15231_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__or2_1
X_09047_ _09047_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _16140_/D sky130_fd_sc_hd__and2_1
XFILLER_0_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold450 hold450/A vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/A vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold483 hold483/A vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 hold494/A vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout930 hold735/X vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__clkbuf_16
Xfanout941 hold129/X vssd1 vssd1 vccd1 vccd1 _14866_/A sky130_fd_sc_hd__buf_6
X_09949_ hold3957/X _10001_/B _09948_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09949_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12987_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _17496_/D sky130_fd_sc_hd__and2_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 input67/X vssd1 vssd1 vccd1 vccd1 hold1150/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 _18096_/Q vssd1 vssd1 vccd1 vccd1 hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ hold3230/X _12302_/B _11910_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _11911_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _16258_/Q vssd1 vssd1 vccd1 vccd1 hold1172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 _17762_/Q vssd1 vssd1 vccd1 vccd1 hold1183/X sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _12918_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _17473_/D sky130_fd_sc_hd__and2_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _08134_/X vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15185_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__or2_1
X_11842_ hold4727/X _12320_/B _11841_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11842_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ hold756/X _14557_/Y _14560_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 hold757/A
+ sky130_fd_sc_hd__o211a_1
X_11773_ _12331_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11773_/Y sky130_fd_sc_hd__nor2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13713_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__or2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _17751_/CLK _16300_/D vssd1 vssd1 vccd1 vccd1 _16300_/Q sky130_fd_sc_hd__dfxtp_1
X_17280_ _17283_/CLK _17280_/D vssd1 vssd1 vccd1 vccd1 _17280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ hold2046/X hold5260/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__mux2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ hold5969/X _14487_/B hold574/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 hold575/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16231_ _17435_/CLK _16231_/D vssd1 vssd1 vccd1 vccd1 _16231_/Q sky130_fd_sc_hd__dfxtp_1
X_13443_ _13737_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10655_ hold1652/X _16709_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16162_ _18013_/CLK _16162_/D vssd1 vssd1 vccd1 vccd1 _16162_/Q sky130_fd_sc_hd__dfxtp_1
X_13374_ _13788_/A _13374_/B vssd1 vssd1 vccd1 vccd1 _13374_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10586_ _10586_/A _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ _15547_/A _15113_/B vssd1 vssd1 vccd1 vccd1 _15113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12325_ _12331_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__nor2_1
X_16093_ _18417_/CLK _16093_/D vssd1 vssd1 vccd1 vccd1 _16093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15044_ _15044_/A hold130/X vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__and2_1
X_12256_ hold5068/X _12347_/B _12255_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _12256_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11207_ _16893_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11207_/X sky130_fd_sc_hd__and3_1
XFILLER_0_142_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12187_ hold4661/X _12377_/B _12186_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ _18073_/Q hold3477/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__mux2_1
X_16995_ _17904_/CLK _16995_/D vssd1 vssd1 vccd1 vccd1 _16995_/Q sky130_fd_sc_hd__dfxtp_1
X_15946_ _17284_/CLK _15946_/D vssd1 vssd1 vccd1 vccd1 hold511/A sky130_fd_sc_hd__dfxtp_1
X_11069_ hold2705/X _16847_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _17715_/CLK _15877_/D vssd1 vssd1 vccd1 vccd1 _15877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17616_ _17739_/CLK _17616_/D vssd1 vssd1 vccd1 vccd1 _17616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ _15221_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__nand2_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ _18392_/CLK _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
X_14759_ hold2746/X _14774_/B _14758_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08280_ _15559_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/X sky130_fd_sc_hd__or2_1
X_17478_ _17480_/CLK _17478_/D vssd1 vssd1 vccd1 vccd1 _17478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_315_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17722_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16429_ _18378_/CLK _16429_/D vssd1 vssd1 vccd1 vccd1 _16429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5405 _16492_/Q vssd1 vssd1 vccd1 vccd1 hold5405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5416 _09829_/X vssd1 vssd1 vccd1 vccd1 _16433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5427 _16476_/Q vssd1 vssd1 vccd1 vccd1 hold5427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5438 _09718_/X vssd1 vssd1 vccd1 vccd1 _16396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4704 _17169_/Q vssd1 vssd1 vccd1 vccd1 hold4704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5449 _11209_/Y vssd1 vssd1 vccd1 vccd1 _16893_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4715 _10507_/X vssd1 vssd1 vccd1 vccd1 _16659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4726 _11455_/X vssd1 vssd1 vccd1 vccd1 _16975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4737 _17218_/Q vssd1 vssd1 vccd1 vccd1 hold4737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4748 _13777_/X vssd1 vssd1 vccd1 vccd1 _17712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4759 _16625_/Q vssd1 vssd1 vccd1 vccd1 hold4759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 _11792_/B vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__buf_4
Xfanout215 _10022_/B vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__buf_4
Xfanout226 _10465_/A2 vssd1 vssd1 vccd1 vccd1 _10568_/B sky130_fd_sc_hd__buf_4
Xfanout237 _09952_/A2 vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__buf_2
X_09803_ hold2000/X _16425_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__mux2_1
Xfanout248 _09494_/X vssd1 vssd1 vccd1 vccd1 _09517_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ hold944/X _08045_/B vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__or2_1
Xfanout259 _12285_/A vssd1 vssd1 vccd1 vccd1 _13794_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ hold362/X _16402_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09665_ hold2532/X _16379_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08616_ _15284_/A _08616_/B vssd1 vssd1 vccd1 vccd1 _15930_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ hold2439/X hold5655/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__mux2_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _09063_/A _08547_/B vssd1 vssd1 vccd1 vccd1 _15897_/D sky130_fd_sc_hd__and2_1
XFILLER_0_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08478_ hold735/X _08500_/B vssd1 vssd1 vccd1 vccd1 _08478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ _10542_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10371_ _10557_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12110_ hold1816/X hold4343/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__mux2_1
Xhold5950 _15866_/Q vssd1 vssd1 vccd1 vccd1 hold5950/X sky130_fd_sc_hd__dlygate4sd3_1
X_13090_ _17562_/Q _17096_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5961 _17868_/Q vssd1 vssd1 vccd1 vccd1 hold5961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5972 data_in[9] vssd1 vssd1 vccd1 vccd1 hold440/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5983 hold6008/X vssd1 vssd1 vccd1 vccd1 hold5983/X sky130_fd_sc_hd__clkbuf_2
Xhold5994 data_in[18] vssd1 vssd1 vccd1 vccd1 hold544/A sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ hold1903/X _17171_/Q _12329_/C vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__mux2_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold38/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout760 _14402_/C1 vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__buf_4
Xfanout771 _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__buf_4
X_15800_ _17731_/CLK _15800_/D vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout782 _14388_/A vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__buf_4
X_13992_ _15553_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__or2_1
X_16780_ _18461_/CLK _16780_/D vssd1 vssd1 vccd1 vccd1 _16780_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout793 fanout816/X vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _17740_/CLK _15731_/D vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfxtp_1
X_12943_ hold2826/X hold3380/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__mux2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18450_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 hold770/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15662_ _17897_/CLK _15662_/D vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ hold2542/X _17469_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux2_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_131 _15207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _18454_/CLK _17401_/D vssd1 vssd1 vccd1 vccd1 _17401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ hold2840/X hold3950/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__mux2_1
X_14613_ hold2403/X _14612_/B _14612_/Y _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14613_/X
+ sky130_fd_sc_hd__o211a_1
X_18381_ _18381_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
X_15593_ _17583_/CLK _15593_/D vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17522_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _17332_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ hold743/X _14541_/B _14543_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 hold744/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _17076_/Q _11762_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _11756_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _11097_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__or2_1
X_17263_ _17263_/CLK _17263_/D vssd1 vssd1 vccd1 vccd1 _17263_/Q sky130_fd_sc_hd__dfxtp_1
X_14475_ _14529_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14475_/X sky130_fd_sc_hd__or2_1
X_11687_ hold2050/X _17053_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16214_ _17691_/CLK _16214_/D vssd1 vssd1 vccd1 vccd1 _16214_/Q sky130_fd_sc_hd__dfxtp_1
X_13426_ hold4805/X _13805_/B _13425_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13426_/X
+ sky130_fd_sc_hd__o211a_1
X_10638_ hold3684/X _10542_/A _10637_/X vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__a21oi_1
X_17194_ _18445_/CLK _17194_/D vssd1 vssd1 vccd1 vccd1 _17194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ _17340_/CLK _16145_/D vssd1 vssd1 vccd1 vccd1 hold713/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13357_ hold4480/X _13856_/B _13356_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ hold3188/X _10560_/A _10568_/X vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _17260_/Q _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__and3_1
X_16076_ _17284_/CLK _16076_/D vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__dfxtp_1
X_13288_ _13281_/X _13287_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__o21a_1
X_15027_ _15189_/A hold2942/X hold302/X vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__mux2_1
X_12239_ hold2072/X hold3368/X _12341_/C vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__mux2_1
Xhold2609 _17867_/Q vssd1 vssd1 vccd1 vccd1 hold2609/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1908 _09147_/X vssd1 vssd1 vccd1 vccd1 _16186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1919 _17777_/Q vssd1 vssd1 vccd1 vccd1 hold1919/X sky130_fd_sc_hd__dlygate4sd3_1
X_07780_ hold173/X vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__inv_2
X_16978_ _17889_/CLK _16978_/D vssd1 vssd1 vccd1 vccd1 _16978_/Q sky130_fd_sc_hd__dfxtp_1
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15929_ _17531_/CLK _15929_/D vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09450_ _09456_/C _09456_/D _09481_/B vssd1 vssd1 vccd1 vccd1 _09450_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08401_ _15515_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
X_09381_ hold521/X _09386_/A _15486_/B1 hold537/X vssd1 vssd1 vccd1 vccd1 _09381_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08332_ hold2464/X _08323_/B _08331_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _08332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08263_ hold2008/X _08262_/B _08262_/Y _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ hold2791/X _08213_/B _08193_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5202 _13567_/X vssd1 vssd1 vccd1 vccd1 _17642_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5213 _17620_/Q vssd1 vssd1 vccd1 vccd1 hold5213/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5224 _16334_/Q vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5235 _11755_/Y vssd1 vssd1 vccd1 vccd1 _17075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4501 _13627_/X vssd1 vssd1 vccd1 vccd1 _17662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5246 _11190_/Y vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4512 _16683_/Q vssd1 vssd1 vccd1 vccd1 hold4512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5257 _16332_/Q vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4523 _09553_/X vssd1 vssd1 vccd1 vccd1 _16341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5268 _11215_/Y vssd1 vssd1 vccd1 vccd1 _16895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5279 _12339_/Y vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4534 _16988_/Q vssd1 vssd1 vccd1 vccd1 hold4534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4545 _13884_/Y vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3800 _11781_/Y vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3811 _17097_/Q vssd1 vssd1 vccd1 vccd1 hold3811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4556 _11425_/X vssd1 vssd1 vccd1 vccd1 _16965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3822 _17583_/Q vssd1 vssd1 vccd1 vccd1 hold3822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4567 _17739_/Q vssd1 vssd1 vccd1 vccd1 hold4567/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3833 _16459_/Q vssd1 vssd1 vccd1 vccd1 hold3833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4578 _15403_/X vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3844 hold5826/X vssd1 vssd1 vccd1 vccd1 hold3844/X sky130_fd_sc_hd__clkbuf_4
Xhold4589 _17616_/Q vssd1 vssd1 vccd1 vccd1 hold4589/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3855 _16455_/Q vssd1 vssd1 vccd1 vccd1 hold3855/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3866 _13806_/Y vssd1 vssd1 vccd1 vccd1 _13807_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3877 _17111_/Q vssd1 vssd1 vccd1 vccd1 hold3877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3888 _16430_/Q vssd1 vssd1 vccd1 vccd1 hold3888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3899 _12358_/Y vssd1 vssd1 vccd1 vccd1 _17276_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _15547_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _09933_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__or2_1
X_09648_ _09951_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__or2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_237_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17749_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10380_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09579_/X sky130_fd_sc_hd__or2_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ _12246_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_0__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_4_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ hold2413/X _12589_/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _11637_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _14529_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__or2_1
X_11472_ _11670_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__or2_1
X_13211_ _13210_/X _16919_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__mux2_1
X_10423_ hold3234/X _10637_/B _10422_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
X_14191_ hold1750/X _14202_/B _14190_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _14191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _13142_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__or2_1
X_10354_ hold4381/X _10640_/B _10353_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10354_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5780 output86/X vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_12
X_13073_ _13073_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__and2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17950_ _18305_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5791 hold5925/X vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__buf_1
X_10285_ hold3453/X _10465_/A2 _10284_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _10285_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12024_ _13794_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__or2_1
X_16901_ _17877_/CLK _16901_/D vssd1 vssd1 vccd1 vccd1 _16901_/Q sky130_fd_sc_hd__dfxtp_1
X_17881_ _17882_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_1
X_16832_ _18035_/CLK _16832_/D vssd1 vssd1 vccd1 vccd1 _16832_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout590 _13049_/Y vssd1 vssd1 vccd1 vccd1 _13311_/C1 sky130_fd_sc_hd__buf_8
XFILLER_0_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ _18054_/CLK _16763_/D vssd1 vssd1 vccd1 vccd1 _16763_/Q sky130_fd_sc_hd__dfxtp_1
X_13975_ hold1744/X _13986_/B _13974_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _13975_/X
+ sky130_fd_sc_hd__o211a_1
X_15714_ _17282_/CLK _15714_/D vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12926_ hold3301/X _12925_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__mux2_1
X_16694_ _18216_/CLK _16694_/D vssd1 vssd1 vccd1 vccd1 _16694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18433_ _18441_/CLK hold946/X vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
X_15645_ _17221_/CLK _15645_/D vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12857_ hold3303/X _12856_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18388_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
X_11808_ _13797_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12788_ hold3052/X _12787_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__mux2_1
X_15576_ _17263_/CLK _15576_/D vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _18421_/CLK _17315_/D vssd1 vssd1 vccd1 vccd1 hold338/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ hold3702/X _11652_/A _11738_/X vssd1 vssd1 vccd1 vccd1 _11739_/Y sky130_fd_sc_hd__a21oi_1
X_14527_ _15099_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ _18385_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _17266_/CLK _17246_/D vssd1 vssd1 vccd1 vccd1 _17246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ hold1569/X _14481_/B _14457_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14458_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13409_ hold2088/X _17590_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__mux2_1
X_17177_ _17583_/CLK _17177_/D vssd1 vssd1 vccd1 vccd1 _17177_/Q sky130_fd_sc_hd__dfxtp_1
X_14389_ _15231_/A hold2709/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _16128_/CLK _16128_/D vssd1 vssd1 vccd1 vccd1 hold525/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _08970_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__and2_1
Xhold3107 _17367_/Q vssd1 vssd1 vccd1 vccd1 hold3107/X sky130_fd_sc_hd__dlygate4sd3_1
X_16059_ _17313_/CLK _16059_/D vssd1 vssd1 vccd1 vccd1 hold576/A sky130_fd_sc_hd__dfxtp_1
Xhold3118 _09394_/X vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3129 _16721_/Q vssd1 vssd1 vccd1 vccd1 hold3129/X sky130_fd_sc_hd__dlygate4sd3_1
X_07901_ hold1273/X _07918_/B _07900_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2406 _14611_/X vssd1 vssd1 vccd1 vccd1 _18099_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08881_ _12428_/A hold256/X vssd1 vssd1 vccd1 vccd1 _16058_/D sky130_fd_sc_hd__and2_1
Xhold2417 _17790_/Q vssd1 vssd1 vccd1 vccd1 hold2417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2428 _14335_/X vssd1 vssd1 vccd1 vccd1 _17967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2439 _18269_/Q vssd1 vssd1 vccd1 vccd1 hold2439/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1705 _14261_/X vssd1 vssd1 vccd1 vccd1 _17931_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ hold2334/X _07865_/B _07831_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _07832_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1716 _15841_/Q vssd1 vssd1 vccd1 vccd1 hold1716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1727 _18061_/Q vssd1 vssd1 vccd1 vccd1 hold1727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 _15753_/Q vssd1 vssd1 vccd1 vccd1 hold1738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 _14476_/X vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09502_ hold5655/X _09998_/B _09501_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09502_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _07804_/A _09477_/A _15314_/A hold629/X vssd1 vssd1 vccd1 vccd1 hold630/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09364_ _09400_/A _09364_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09364_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08315_ _15539_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08315_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _15517_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__or2_1
XANTENNA_31 _17524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _14986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_53 _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _15525_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_64 hold335/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_75 hold800/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_86 hold5845/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_97 _14545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ hold756/X _08225_/B vssd1 vssd1 vccd1 vccd1 _08177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5010 _09667_/X vssd1 vssd1 vccd1 vccd1 _16379_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5021 _17232_/Q vssd1 vssd1 vccd1 vccd1 hold5021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5032 _16590_/Q vssd1 vssd1 vccd1 vccd1 hold5032/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5043 _11833_/X vssd1 vssd1 vccd1 vccd1 _17101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5054 _16005_/Q vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5065 _11317_/X vssd1 vssd1 vccd1 vccd1 _16929_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4320 _09706_/X vssd1 vssd1 vccd1 vccd1 _16392_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5076 _16506_/Q vssd1 vssd1 vccd1 vccd1 hold5076/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4331 _17725_/Q vssd1 vssd1 vccd1 vccd1 hold4331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5087 _13366_/X vssd1 vssd1 vccd1 vccd1 _17575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4342 _10756_/X vssd1 vssd1 vccd1 vccd1 _16742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5098 _16451_/Q vssd1 vssd1 vccd1 vccd1 hold5098/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4353 _16801_/Q vssd1 vssd1 vccd1 vccd1 hold4353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4364 _11029_/X vssd1 vssd1 vccd1 vccd1 _16833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3630 _16542_/Q vssd1 vssd1 vccd1 vccd1 hold3630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4375 _16580_/Q vssd1 vssd1 vccd1 vccd1 hold4375/X sky130_fd_sc_hd__dlygate4sd3_1
X_10070_ _16514_/Q _10070_/B _10271_/S vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__and3_1
Xhold3641 _10627_/Y vssd1 vssd1 vccd1 vccd1 _16699_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4386 _13540_/X vssd1 vssd1 vccd1 vccd1 _17633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3652 _13827_/Y vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4397 _16992_/Q vssd1 vssd1 vccd1 vccd1 hold4397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3663 _10572_/Y vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3674 _10576_/Y vssd1 vssd1 vccd1 vccd1 _16682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2940 _17926_/Q vssd1 vssd1 vccd1 vccd1 hold2940/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3685 _10638_/Y vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3696 _16720_/Q vssd1 vssd1 vccd1 vccd1 hold3696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2951 _16266_/Q vssd1 vssd1 vccd1 vccd1 hold2951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2962 _08400_/X vssd1 vssd1 vccd1 vccd1 _15830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 _18110_/Q vssd1 vssd1 vccd1 vccd1 hold2973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2984 _14925_/X vssd1 vssd1 vccd1 vccd1 _18249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2995 _18190_/Q vssd1 vssd1 vccd1 vccd1 hold2995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ hold2648/X _17707_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__mux2_1
X_10972_ hold5572/X _09992_/B _10971_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _12777_/A _12711_/B vssd1 vssd1 vccd1 vccd1 _17413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13691_ hold1501/X _17684_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13692_/B sky130_fd_sc_hd__mux2_1
X_15430_ hold200/X _09365_/B _09362_/D hold374/X _15428_/X vssd1 vssd1 vccd1 vccd1
+ _15432_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12642_ _12885_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _17390_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _16300_/Q _09362_/A _09392_/B hold515/X _15360_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/D sky130_fd_sc_hd__a221o_1
X_12573_ _12996_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _17367_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17100_ _17253_/CLK _17100_/D vssd1 vssd1 vccd1 vccd1 _17100_/Q sky130_fd_sc_hd__dfxtp_1
X_11524_ hold4881/X _12305_/B _11523_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11524_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _15207_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__or2_1
X_15292_ _15489_/A _15292_/B _15292_/C _15292_/D vssd1 vssd1 vccd1 vccd1 _15292_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18080_ _18080_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17031_ _17879_/CLK _17031_/D vssd1 vssd1 vccd1 vccd1 _17031_/Q sky130_fd_sc_hd__dfxtp_1
X_14243_ hold1144/X _14266_/B _14242_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14243_/X
+ sky130_fd_sc_hd__o211a_1
X_11455_ hold4725/X _12323_/B _11454_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ hold1996/X _16626_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__mux2_1
X_14174_ _15193_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14174_/X sky130_fd_sc_hd__or2_1
X_11386_ hold4514/X _11798_/B _11385_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11386_/X
+ sky130_fd_sc_hd__o211a_1
X_13125_ _13124_/X hold3633/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__mux2_1
X_10337_ hold2797/X hold4030/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__mux2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _17523_/Q _17522_/Q _13056_/C _13056_/D vssd1 vssd1 vccd1 vccd1 _13056_/X
+ sky130_fd_sc_hd__and4b_4
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _18061_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
X_10268_ hold3029/X _16580_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10269_/B sky130_fd_sc_hd__mux2_1
X_12007_ hold3340/X _12302_/B _12006_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _17896_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
X_10199_ hold2139/X hold3210/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_159_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18230_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16815_ _18050_/CLK _16815_/D vssd1 vssd1 vccd1 vccd1 _16815_/Q sky130_fd_sc_hd__dfxtp_1
X_17795_ _17827_/CLK hold870/X vssd1 vssd1 vccd1 vccd1 hold869/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16746_ _18042_/CLK _16746_/D vssd1 vssd1 vccd1 vccd1 _16746_/Q sky130_fd_sc_hd__dfxtp_1
X_13958_ hold826/X _13992_/B vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ _12909_/A _12909_/B vssd1 vssd1 vccd1 vccd1 _17479_/D sky130_fd_sc_hd__and2_1
X_16677_ _18267_/CLK _16677_/D vssd1 vssd1 vccd1 vccd1 _16677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ _07786_/Y _16286_/Q hold927/X _10763_/S vssd1 vssd1 vccd1 vccd1 hold928/A
+ sky130_fd_sc_hd__a31oi_1
X_18416_ _18416_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15628_ _17724_/CLK _15628_/D vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ _18373_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08100_ _14786_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09080_ _14980_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _18420_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08031_ _15545_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 input40/A vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_17229_ _17718_/CLK _17229_/D vssd1 vssd1 vccd1 vccd1 _17229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput51 input51/A vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_6
Xhold802 hold802/A vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 hold813/A vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold824 hold857/X vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 hold835/A vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 la_data_in[5] vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _13062_/A _10022_/B _09981_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _09982_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold879 input52/X vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ _12402_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _16084_/D sky130_fd_sc_hd__and2_1
Xhold2203 _18119_/Q vssd1 vssd1 vccd1 vccd1 hold2203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 _12679_/X vssd1 vssd1 vccd1 vccd1 hold2214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2225 _12647_/X vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2236 _17855_/Q vssd1 vssd1 vccd1 vccd1 hold2236/X sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ hold14/X _16051_/Q _08864_/S vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__mux2_1
Xhold1502 _08261_/X vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2247 _14490_/X vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 _18340_/Q vssd1 vssd1 vccd1 vccd1 hold2258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _15852_/Q vssd1 vssd1 vccd1 vccd1 hold1513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 _15080_/X vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 _14721_/X vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 hold5822/X vssd1 vssd1 vccd1 vccd1 _13043_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ hold949/X _14980_/A _15519_/A _15517_/A vssd1 vssd1 vccd1 vccd1 _07817_/C
+ sky130_fd_sc_hd__or4_1
Xhold1546 _18000_/Q vssd1 vssd1 vccd1 vccd1 hold1546/X sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ _13056_/C _13030_/A vssd1 vssd1 vccd1 vccd1 _13046_/D sky130_fd_sc_hd__nand2_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 _18160_/Q vssd1 vssd1 vccd1 vccd1 hold1557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1568 _15092_/X vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 _09419_/X vssd1 vssd1 vccd1 vccd1 _16295_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09416_ _09438_/B _16294_/Q vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09347_ _09400_/A _09363_/B _09351_/B vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _12813_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _16250_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08229_ _08504_/A hold607/X vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__or2_4
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11240_ hold1365/X hold3778/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11241_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _16881_/Q _11171_/B _11171_/C vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4150 _11134_/X vssd1 vssd1 vccd1 vccd1 _16868_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10122_ _10506_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10122_/X sky130_fd_sc_hd__or2_1
Xhold4161 _17623_/Q vssd1 vssd1 vccd1 vccd1 hold4161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4172 _17158_/Q vssd1 vssd1 vccd1 vccd1 hold4172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4183 _10360_/X vssd1 vssd1 vccd1 vccd1 _16610_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4194 _16657_/Q vssd1 vssd1 vccd1 vccd1 hold4194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3460 _09397_/X vssd1 vssd1 vccd1 vccd1 _16285_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14930_ _15199_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14930_/X sky130_fd_sc_hd__or2_1
X_10053_ _13254_/A _09975_/A _10052_/X vssd1 vssd1 vccd1 vccd1 _10053_/Y sky130_fd_sc_hd__a21oi_1
Xhold3471 _12046_/X vssd1 vssd1 vccd1 vccd1 _17172_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3482 _17736_/Q vssd1 vssd1 vccd1 vccd1 hold3482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3493 _17445_/Q vssd1 vssd1 vccd1 vccd1 hold3493/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_252_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17736_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2770 _13961_/X vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14861_ hold2736/X _14880_/B _14860_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14861_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2781 _15854_/Q vssd1 vssd1 vccd1 vccd1 hold2781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2792 _08194_/X vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16600_ _18190_/CLK _16600_/D vssd1 vssd1 vccd1 vccd1 _16600_/Q sky130_fd_sc_hd__dfxtp_1
X_13812_ hold3883/X _13716_/A _13811_/X vssd1 vssd1 vccd1 vccd1 _13812_/Y sky130_fd_sc_hd__a21oi_1
X_17580_ _17740_/CLK _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
X_14792_ _15185_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14792_/X sky130_fd_sc_hd__or2_1
X_16531_ _18217_/CLK _16531_/D vssd1 vssd1 vccd1 vccd1 _16531_/Q sky130_fd_sc_hd__dfxtp_1
X_13743_ _13776_/A _13743_/B vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__or2_1
X_10955_ hold2161/X _16809_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16462_ _18416_/CLK _16462_/D vssd1 vssd1 vccd1 vccd1 _16462_/Q sky130_fd_sc_hd__dfxtp_1
X_13674_ _13674_/A _13674_/B vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__or2_1
X_10886_ hold422/X hold5417/X _11753_/C vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18201_ _18230_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
X_15413_ _15490_/A1 _15405_/X _15412_/X _15490_/B1 _18417_/Q vssd1 vssd1 vccd1 vccd1
+ _15413_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ hold1313/X _17386_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16393_ _18339_/CLK _16393_/D vssd1 vssd1 vccd1 vccd1 _16393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18132_ _18222_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ _15344_/A _15344_/B vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__and2_1
X_12556_ hold1112/X _17363_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11507_ hold1253/X _16993_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__mux2_1
X_18063_ _18063_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
X_15275_ _15275_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__or2_1
X_12487_ hold5/X _08598_/B _08999_/B _12486_/X _15414_/A vssd1 vssd1 vccd1 vccd1 hold6/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold109 hold13/X vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _17798_/CLK _17014_/D vssd1 vssd1 vccd1 vccd1 _17014_/Q sky130_fd_sc_hd__dfxtp_1
X_11438_ hold1383/X _16970_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__mux2_1
X_14226_ _15517_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14226_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14157_ hold969/X _14148_/B _14156_/X _15504_/A vssd1 vssd1 vccd1 vccd1 hold970/A
+ sky130_fd_sc_hd__o211a_1
X_11369_ hold869/X _16947_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ hold3616/X _13107_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__mux2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _15541_/A _14094_/B vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__nand2_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13039_/A _13039_/B vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__and2_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _18042_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_1
X_17847_ _17880_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08580_ hold251/X hold390/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__mux2_1
X_17778_ _17905_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _18033_/CLK _16729_/D vssd1 vssd1 vccd1 vccd1 _16729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ hold1950/X _09218_/B _09200_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09201_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17487_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09132_ _15515_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _16148_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08014_ hold2626/X _08029_/B _08013_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _08014_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 hold610/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 la_data_in[26] vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 hold643/A vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 input61/X vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold665 hold665/A vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 hold676/A vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold687 hold687/A vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 hold698/A vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ hold2693/X _16479_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__mux2_1
Xhold2000 _18338_/Q vssd1 vssd1 vccd1 vccd1 hold2000/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2011 _07919_/X vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2022 _18201_/Q vssd1 vssd1 vccd1 vccd1 hold2022/X sky130_fd_sc_hd__dlygate4sd3_1
X_08916_ hold149/X hold458/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__mux2_1
Xhold2033 _08210_/X vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 _15629_/Q vssd1 vssd1 vccd1 vccd1 hold2044/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _18369_/Q hold5496/X _11066_/S vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__mux2_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _14125_/X vssd1 vssd1 vccd1 vccd1 _17866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2055 _14107_/X vssd1 vssd1 vccd1 vccd1 _17858_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _14189_/X vssd1 vssd1 vccd1 vccd1 _17897_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2066 _17852_/Q vssd1 vssd1 vccd1 vccd1 hold2066/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1332 _18346_/Q vssd1 vssd1 vccd1 vccd1 hold1332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2077 _07907_/X vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _15196_/X vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _15364_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _16042_/D sky130_fd_sc_hd__and2_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2088 _15879_/Q vssd1 vssd1 vccd1 vccd1 hold2088/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1354 _14099_/X vssd1 vssd1 vccd1 vccd1 _17854_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2099 _15164_/X vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1365 _18430_/Q vssd1 vssd1 vccd1 vccd1 hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1376 _07971_/X vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ _15482_/A hold150/X vssd1 vssd1 vccd1 vccd1 _16009_/D sky130_fd_sc_hd__and2_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 _15777_/Q vssd1 vssd1 vccd1 vccd1 hold1387/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _08473_/X vssd1 vssd1 vccd1 vccd1 _15865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _11031_/A _10740_/B vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ _11136_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12410_ _12426_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _17298_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ hold4955/X _13847_/B _13389_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13390_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12341_ _17271_/Q _12341_/B _12341_/C vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__and3_1
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15060_ _15060_/A hold363/X vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ hold2109/X _17248_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__mux2_1
X_14011_ hold993/X _14036_/B _14010_/X _13943_/A vssd1 vssd1 vccd1 vccd1 hold994/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ hold5318/X _11031_/A _11222_/X vssd1 vssd1 vccd1 vccd1 _11223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ hold5294/X _11136_/A _11153_/X vssd1 vssd1 vccd1 vccd1 _11154_/Y sky130_fd_sc_hd__a21oi_1
X_10105_ hold3210/X _10649_/B _10104_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10105_/X
+ sky130_fd_sc_hd__o211a_1
X_15962_ _18425_/CLK _15962_/D vssd1 vssd1 vccd1 vccd1 hold614/A sky130_fd_sc_hd__dfxtp_1
X_11085_ _11097_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17701_ _17701_/CLK _17701_/D vssd1 vssd1 vccd1 vccd1 _17701_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3290 _12866_/X vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14913_ _14913_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14962_/B sky130_fd_sc_hd__or2_4
X_10036_ _11194_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__nor2_1
X_15893_ _17343_/CLK _15893_/D vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__dfxtp_1
X_17632_ _17731_/CLK _17632_/D vssd1 vssd1 vccd1 vccd1 _17632_/Q sky130_fd_sc_hd__dfxtp_1
X_14844_ _15129_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ _17723_/CLK _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
X_14775_ hold2191/X _14774_/B _14774_/Y _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14775_/X
+ sky130_fd_sc_hd__o211a_1
X_11987_ hold2860/X _17153_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__mux2_1
X_16514_ _18395_/CLK _16514_/D vssd1 vssd1 vccd1 vccd1 _16514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13726_ hold4207/X _13829_/B _13725_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13726_/X
+ sky130_fd_sc_hd__o211a_1
X_10938_ _11670_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__or2_1
X_17494_ _17494_/CLK _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16445_ _18358_/CLK _16445_/D vssd1 vssd1 vccd1 vccd1 _16445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13657_ hold3570/X _13847_/B _13656_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13657_/X
+ sky130_fd_sc_hd__o211a_1
X_10869_ _11061_/A _10869_/B vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__or2_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ hold3253/X _12607_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__mux2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _18353_/CLK _16376_/D vssd1 vssd1 vccd1 vccd1 _16376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ hold3573/X _13886_/B _13587_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13588_/X
+ sky130_fd_sc_hd__o211a_1
X_18115_ _18266_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
X_15327_ hold375/X _09357_/A _15484_/B1 hold322/X _15326_/X vssd1 vssd1 vccd1 vccd1
+ _15332_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_136_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12539_ hold3586/X _12538_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5609 _10969_/X vssd1 vssd1 vccd1 vccd1 _16813_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ _18046_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
X_15258_ hold460/X _15484_/A2 _15451_/A2 _17286_/Q vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4908 _13327_/X vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4919 _17153_/Q vssd1 vssd1 vccd1 vccd1 hold4919/X sky130_fd_sc_hd__dlygate4sd3_1
X_14209_ hold1977/X _14202_/B _14208_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14209_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15189_ _15189_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_174_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18067_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout408 _14286_/Y vssd1 vssd1 vccd1 vccd1 _14326_/B sky130_fd_sc_hd__buf_4
Xfanout419 _14105_/A2 vssd1 vssd1 vccd1 vccd1 _14094_/B sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_103_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17342_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09750_ _09954_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__or2_1
X_08701_ hold219/X hold723/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__mux2_1
X_09681_ _10491_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08632_ _12430_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _15938_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _09063_/A hold182/X vssd1 vssd1 vccd1 vccd1 _15905_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08494_ _14726_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09115_ hold2697/X _09119_/A2 _09114_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _09115_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ hold149/X hold287/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09047_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold440 hold440/A vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold451/A vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold473 hold473/A vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout920 hold730/X vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__buf_12
Xfanout931 hold735/X vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__clkbuf_16
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__or2_1
Xfanout942 hold747/X vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__buf_12
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _09975_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__or2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 _16150_/Q vssd1 vssd1 vccd1 vccd1 hold1140/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _08302_/X vssd1 vssd1 vccd1 vccd1 _15784_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _14605_/X vssd1 vssd1 vccd1 vccd1 _18096_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _12210_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__or2_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1173 _09296_/X vssd1 vssd1 vccd1 vccd1 _16258_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ hold3259/X _12889_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__mux2_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _13908_/X vssd1 vssd1 vccd1 vccd1 _13909_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _18029_/Q vssd1 vssd1 vccd1 vccd1 hold1195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _12093_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__or2_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ hold5236/X _12051_/A _11771_/X vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _15492_/A _14573_/B _18075_/Q vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__a21o_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ hold1087/X _17624_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ hold4035/X _11201_/B _10722_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _10723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ hold573/X _14499_/B vssd1 vssd1 vccd1 vccd1 hold574/A sky130_fd_sc_hd__or2_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _17439_/CLK _16230_/D vssd1 vssd1 vccd1 vccd1 _16230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ hold1864/X hold4281/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__mux2_1
X_10654_ hold3202/X _11171_/B _10653_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _10654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ hold1700/X hold4169/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__mux2_1
X_16161_ _18013_/CLK _16161_/D vssd1 vssd1 vccd1 vccd1 _16161_/Q sky130_fd_sc_hd__dfxtp_1
X_10585_ _10588_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15112_ hold2258/X _15113_/B _15111_/Y _15050_/A vssd1 vssd1 vccd1 vccd1 _15112_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12324_ hold3835/X _12036_/A _12323_/X vssd1 vssd1 vccd1 vccd1 _12324_/Y sky130_fd_sc_hd__a21oi_1
X_16092_ _18413_/CLK _16092_/D vssd1 vssd1 vccd1 vccd1 hold552/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _12255_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12255_/X sky130_fd_sc_hd__or2_1
X_15043_ hold129/X _18307_/Q hold302/A vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ _12331_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _11206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12186_ _12282_/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__or2_1
X_11137_ hold5590/X _11156_/B _11136_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _11137_/X
+ sky130_fd_sc_hd__o211a_1
X_16994_ _17905_/CLK _16994_/D vssd1 vssd1 vccd1 vccd1 _16994_/Q sky130_fd_sc_hd__dfxtp_1
X_15945_ _17292_/CLK _15945_/D vssd1 vssd1 vccd1 vccd1 hold382/A sky130_fd_sc_hd__dfxtp_1
X_11068_ hold5703/X _09992_/B _11067_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _11068_/X
+ sky130_fd_sc_hd__o211a_1
X_10019_ _16497_/Q _10025_/B _10025_/C vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__and3_1
X_15876_ _17737_/CLK _15876_/D vssd1 vssd1 vccd1 vccd1 _15876_/Q sky130_fd_sc_hd__dfxtp_1
X_17615_ _17647_/CLK _17615_/D vssd1 vssd1 vccd1 vccd1 _17615_/Q sky130_fd_sc_hd__dfxtp_1
X_14827_ hold2875/X _14828_/B _14826_/Y _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14827_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _18392_/CLK _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14758_ _15205_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ hold1509/X hold4333/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17477_ _17480_/CLK _17477_/D vssd1 vssd1 vccd1 vccd1 _17477_/Q sky130_fd_sc_hd__dfxtp_1
X_14689_ hold2955/X _14720_/B _14688_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14689_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ _18334_/CLK _16428_/D vssd1 vssd1 vccd1 vccd1 _16428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16359_ _18304_/CLK _16359_/D vssd1 vssd1 vccd1 vccd1 _16359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5406 _09910_/X vssd1 vssd1 vccd1 vccd1 _16460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5417 _16786_/Q vssd1 vssd1 vccd1 vccd1 hold5417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5428 _09862_/X vssd1 vssd1 vccd1 vccd1 _16444_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5439 _16401_/Q vssd1 vssd1 vccd1 vccd1 hold5439/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4705 _11941_/X vssd1 vssd1 vccd1 vccd1 _17137_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18029_ _18066_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4716 _16793_/Q vssd1 vssd1 vccd1 vccd1 hold4716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4727 _17136_/Q vssd1 vssd1 vccd1 vccd1 hold4727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4738 _12088_/X vssd1 vssd1 vccd1 vccd1 _17186_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4749 _16944_/Q vssd1 vssd1 vccd1 vccd1 hold4749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 fanout209/X vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__buf_4
XFILLER_0_157_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout216 _10022_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__buf_4
X_09802_ hold5496/X _09992_/B _09801_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09802_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout227 _10897_/A2 vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__buf_4
Xfanout238 _10601_/B vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__buf_4
Xfanout249 _13713_/A vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__buf_4
X_07994_ hold816/X _14681_/A vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__or2_4
X_09733_ hold5379/X _10025_/B _09732_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09733_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ hold5017/X _10070_/B _09663_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09664_/X
+ sky130_fd_sc_hd__o211a_1
X_08615_ hold126/X hold415/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__mux2_1
X_09595_ hold5134/X _10073_/B _09594_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09595_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_71_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17289_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ hold47/X hold434/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08547_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08477_ hold1700/X _08486_/B _08476_/X _13753_/C1 vssd1 vssd1 vccd1 vccd1 _08477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ hold1720/X _16614_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _15491_/A hold671/X vssd1 vssd1 vccd1 vccd1 _16131_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5940 hold5997/X vssd1 vssd1 vccd1 vccd1 hold5940/X sky130_fd_sc_hd__buf_1
XFILLER_0_131_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5951 _15840_/Q vssd1 vssd1 vccd1 vccd1 hold5951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5962 _15784_/Q vssd1 vssd1 vccd1 vccd1 hold5962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5973 _17869_/Q vssd1 vssd1 vccd1 vccd1 hold5973/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ hold4865/X _12362_/B _12039_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _12040_/X
+ sky130_fd_sc_hd__o211a_1
Xhold270 hold814/X vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__buf_4
Xhold5984 _18004_/Q vssd1 vssd1 vccd1 vccd1 hold5984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5995 _18412_/Q vssd1 vssd1 vccd1 vccd1 hold5995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__clkbuf_2
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout750 fanout763/X vssd1 vssd1 vccd1 vccd1 _12142_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout761 _14402_/C1 vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__buf_4
Xfanout772 _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__clkbuf_4
X_13991_ hold1428/X _13986_/B _13990_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout783 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout794 _15060_/A vssd1 vssd1 vccd1 vccd1 _15054_/A sky130_fd_sc_hd__buf_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _17732_/CLK _15730_/D vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12951_/A _12942_/B vssd1 vssd1 vccd1 vccd1 _17490_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _17205_/CLK _15661_/D vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _14850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _12885_/A _12873_/B vssd1 vssd1 vccd1 vccd1 _17467_/D sky130_fd_sc_hd__and2_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_132 _13051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _18454_/CLK _17400_/D vssd1 vssd1 vccd1 vccd1 _17400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14774_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__nand2_1
X_18380_ _18380_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11824_ hold3320/X _13811_/B _11823_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _11824_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _17906_/CLK _15592_/D vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17331_ _17331_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _17331_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ hold730/X _14545_/B vssd1 vssd1 vccd1 vccd1 _14543_/X sky130_fd_sc_hd__or2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _12331_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__nor2_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17262_ _17262_/CLK _17262_/D vssd1 vssd1 vccd1 vccd1 _17262_/Q sky130_fd_sc_hd__dfxtp_1
X_10706_ hold2844/X hold3784/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__mux2_1
X_14474_ hold2889/X _14481_/B _14473_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14474_/X
+ sky130_fd_sc_hd__o211a_1
X_11686_ hold5090/X _12323_/B _11685_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11686_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16213_ _17447_/CLK _16213_/D vssd1 vssd1 vccd1 vccd1 _16213_/Q sky130_fd_sc_hd__dfxtp_1
X_13425_ _13710_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _13425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ _16703_/Q _10637_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__and3_1
X_17193_ _17257_/CLK _17193_/D vssd1 vssd1 vccd1 vccd1 _17193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _17343_/CLK _16144_/D vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__dfxtp_1
X_10568_ _16680_/Q _10568_/B _10568_/C vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and3_1
X_13356_ _13770_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _13822_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _17259_/D sky130_fd_sc_hd__nor2_1
X_16075_ _17341_/CLK _16075_/D vssd1 vssd1 vccd1 vccd1 hold688/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10499_ hold1612/X hold4194/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__mux2_1
X_13287_ _13311_/A1 _13285_/X _13286_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13287_/X
+ sky130_fd_sc_hd__o211a_1
X_15026_ _15026_/A _15026_/B vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__and2_1
X_12238_ hold3515/X _12347_/B _12237_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12238_/X
+ sky130_fd_sc_hd__o211a_1
X_12169_ hold5044/X _12347_/B _12168_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _12169_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1909 _18103_/Q vssd1 vssd1 vccd1 vccd1 hold1909/X sky130_fd_sc_hd__dlygate4sd3_1
X_16977_ _17923_/CLK _16977_/D vssd1 vssd1 vccd1 vccd1 _16977_/Q sky130_fd_sc_hd__dfxtp_1
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ _17531_/CLK _15928_/D vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15859_ _17730_/CLK _15859_/D vssd1 vssd1 vccd1 vccd1 _15859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ hold2961/X _08440_/A2 _08399_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _08400_/X
+ sky130_fd_sc_hd__o211a_1
X_09380_ hold597/X _09365_/B _15477_/A2 vssd1 vssd1 vccd1 vccd1 _09383_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08331_ hold800/X _08335_/B vssd1 vssd1 vccd1 vccd1 _08331_/X sky130_fd_sc_hd__or2_1
X_17529_ _17530_/CLK _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _15000_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08193_ _15527_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5203 _17652_/Q vssd1 vssd1 vccd1 vccd1 hold5203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5214 _13405_/X vssd1 vssd1 vccd1 vccd1 _17588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5225 _10011_/Y vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5236 _16921_/Q vssd1 vssd1 vccd1 vccd1 hold5236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4502 _17234_/Q vssd1 vssd1 vccd1 vccd1 hold4502/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5247 _11191_/Y vssd1 vssd1 vccd1 vccd1 _16887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4513 _10483_/X vssd1 vssd1 vccd1 vccd1 _16651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5258 _10005_/Y vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5269 _16339_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4524 _16943_/Q vssd1 vssd1 vccd1 vccd1 hold4524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4535 _11398_/X vssd1 vssd1 vccd1 vccd1 _16956_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4546 _13885_/Y vssd1 vssd1 vccd1 vccd1 _17748_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3801 _11782_/Y vssd1 vssd1 vccd1 vccd1 _17084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4557 _17660_/Q vssd1 vssd1 vccd1 vccd1 hold4557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3812 _12300_/Y vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3823 _13869_/Y vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4568 _13762_/X vssd1 vssd1 vccd1 vccd1 _17707_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3834 _09811_/X vssd1 vssd1 vccd1 vccd1 _16427_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4579 _17016_/Q vssd1 vssd1 vccd1 vccd1 hold4579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3845 _15263_/X vssd1 vssd1 vccd1 vccd1 _15264_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3856 _09799_/X vssd1 vssd1 vccd1 vccd1 _16423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3867 _13807_/Y vssd1 vssd1 vccd1 vccd1 _17722_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3878 _12342_/Y vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3889 _09724_/X vssd1 vssd1 vccd1 vccd1 _16398_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07977_ hold1943/X _07978_/B _07976_/Y _08159_/A vssd1 vssd1 vccd1 vccd1 _07977_/X
+ sky130_fd_sc_hd__o211a_1
X_09716_ hold1670/X _16396_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09717_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ hold2074/X _16373_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__mux2_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09578_ hold847/X _13270_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _12422_/A hold514/X vssd1 vssd1 vccd1 vccd1 _15889_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_277_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ hold2066/X _17004_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_206_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17894_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ hold1941/X _16981_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _10422_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__or2_1
X_13210_ _17577_/Q _17111_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14190_ _14529_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14190_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13141_ _13140_/X hold5901/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
X_10353_ _10554_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5770 output85/X vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_12
X_13072_ _13065_/X _13071_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17527_/D sky130_fd_sc_hd__o21a_1
Xhold5781 hold5920/X vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10284_ _10560_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__or2_1
Xhold5792 hold5792/A vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_12
XFILLER_0_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12023_ hold2295/X hold3474/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__mux2_1
X_16900_ _17844_/CLK _16900_/D vssd1 vssd1 vccd1 vccd1 _16900_/Q sky130_fd_sc_hd__dfxtp_1
X_17880_ _17880_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
X_16831_ _18066_/CLK _16831_/D vssd1 vssd1 vccd1 vccd1 _16831_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout580 _14572_/X vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__buf_6
Xfanout591 _12814_/S vssd1 vssd1 vccd1 vccd1 _12805_/S sky130_fd_sc_hd__clkbuf_8
X_16762_ _18032_/CLK _16762_/D vssd1 vssd1 vccd1 vccd1 _16762_/Q sky130_fd_sc_hd__dfxtp_1
X_13974_ _14529_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13974_/X sky130_fd_sc_hd__or2_1
X_15713_ _17281_/CLK _15713_/D vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ hold1075/X _17486_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__mux2_1
X_16693_ _18219_/CLK _16693_/D vssd1 vssd1 vccd1 vccd1 _16693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18432_ _18432_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
X_15644_ _17844_/CLK _15644_/D vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ hold1619/X _17463_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18363_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
X_11807_ _15718_/Q _17093_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _17232_/CLK _15575_/D vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ hold2624/X _17440_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17314_ _17314_/CLK _17314_/D vssd1 vssd1 vccd1 vccd1 hold536/A sky130_fd_sc_hd__dfxtp_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ hold2848/X _14541_/B _14525_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14526_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18294_ _18358_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _17070_/Q _11747_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17245_ _17743_/CLK _17245_/D vssd1 vssd1 vccd1 vccd1 _17245_/Q sky130_fd_sc_hd__dfxtp_1
X_14457_ _15191_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14457_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ hold804/X _17047_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ hold4931/X _13886_/B _13407_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13408_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17176_ _17208_/CLK _17176_/D vssd1 vssd1 vccd1 vccd1 _17176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14388_ _14388_/A _14388_/B vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16127_ _17531_/CLK _16127_/D vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__dfxtp_1
X_13339_ hold3293/X _13862_/B _13338_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16058_ _17289_/CLK _16058_/D vssd1 vssd1 vccd1 vccd1 _16058_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3108 _12572_/X vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3119 _17442_/Q vssd1 vssd1 vccd1 vccd1 hold3119/X sky130_fd_sc_hd__dlygate4sd3_1
X_15009_ hold775/X _15004_/B _15008_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 hold776/A
+ sky130_fd_sc_hd__o211a_1
X_07900_ _14517_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07900_/X sky130_fd_sc_hd__or2_1
Xhold2407 _18445_/Q vssd1 vssd1 vccd1 vccd1 hold2407/X sky130_fd_sc_hd__dlygate4sd3_1
X_08880_ hold41/X _16058_/Q _08932_/S vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__mux2_1
Xhold2418 _13967_/X vssd1 vssd1 vccd1 vccd1 _17790_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2429 _17941_/Q vssd1 vssd1 vccd1 vccd1 hold2429/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1706 _18188_/Q vssd1 vssd1 vccd1 vccd1 hold1706/X sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ _14218_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07831_/X sky130_fd_sc_hd__or2_1
Xhold1717 _08422_/X vssd1 vssd1 vccd1 vccd1 _15841_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 _14530_/X vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _08237_/X vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09501_ _09903_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__or2_1
XFILLER_0_177_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ hold616/X _16302_/Q vssd1 vssd1 vccd1 vccd1 hold629/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ _09400_/A _09363_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09363_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08314_ hold1992/X _08323_/B _08313_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09294_ hold1646/X _09338_/A2 _09293_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09294_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_10 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_32 _18421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ hold1418/X _08262_/B _08244_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_54 hold892/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_65 hold335/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_76 hold883/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_87 hold5851/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ hold2654/X _08209_/B _08175_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08176_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_98 _14545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5000 _09847_/X vssd1 vssd1 vccd1 vccd1 _16439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5011 _16563_/Q vssd1 vssd1 vccd1 vccd1 hold5011/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5022 _12130_/X vssd1 vssd1 vccd1 vccd1 _17200_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5033 _10204_/X vssd1 vssd1 vccd1 vccd1 _16558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5044 _17245_/Q vssd1 vssd1 vccd1 vccd1 hold5044/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4310 _09865_/X vssd1 vssd1 vccd1 vccd1 _16445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5055 _15363_/X vssd1 vssd1 vccd1 vccd1 _15364_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4321 _16596_/Q vssd1 vssd1 vccd1 vccd1 hold4321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5066 _17640_/Q vssd1 vssd1 vccd1 vccd1 hold5066/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4332 _13720_/X vssd1 vssd1 vccd1 vccd1 _17693_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5077 _09952_/X vssd1 vssd1 vccd1 vccd1 _16474_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4343 _17194_/Q vssd1 vssd1 vccd1 vccd1 hold4343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5088 _17163_/Q vssd1 vssd1 vccd1 vccd1 hold5088/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5099 _09787_/X vssd1 vssd1 vccd1 vccd1 _16419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4354 _10837_/X vssd1 vssd1 vccd1 vccd1 _16769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4365 _16608_/Q vssd1 vssd1 vccd1 vccd1 hold4365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3620 _10617_/Y vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4376 _10174_/X vssd1 vssd1 vccd1 vccd1 _16548_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3631 _10635_/Y vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4387 _16693_/Q vssd1 vssd1 vccd1 vccd1 hold4387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3642 _16545_/Q vssd1 vssd1 vccd1 vccd1 hold3642/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3653 _13828_/Y vssd1 vssd1 vccd1 vccd1 _17729_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4398 _11410_/X vssd1 vssd1 vccd1 vccd1 _16960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3664 _10573_/Y vssd1 vssd1 vccd1 vccd1 _16681_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2930 _18141_/Q vssd1 vssd1 vccd1 vccd1 hold2930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3675 _16350_/Q vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3686 _10639_/Y vssd1 vssd1 vccd1 vccd1 _16703_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2941 _14251_/X vssd1 vssd1 vccd1 vccd1 _17926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3697 _11169_/Y vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2952 _09312_/X vssd1 vssd1 vccd1 vccd1 _16266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 _15615_/Q vssd1 vssd1 vccd1 vccd1 hold2963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2974 _14635_/X vssd1 vssd1 vccd1 vccd1 _18110_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2985 _18027_/Q vssd1 vssd1 vccd1 vccd1 hold2985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2996 _14801_/X vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10971_ _11067_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10971_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ hold3520/X _12709_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__mux2_1
X_13690_ hold5102/X _13883_/B _13689_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13690_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ hold3081/X _12640_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15360_ hold619/X _09367_/A _09392_/A hold716/X vssd1 vssd1 vccd1 vccd1 _15360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ hold3107/X _12571_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14311_ hold2601/X _14333_/A2 _14310_/X _14378_/A vssd1 vssd1 vccd1 vccd1 _14311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ _12018_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__or2_1
X_15291_ _16293_/Q _15477_/A2 _15487_/B1 hold482/X _15290_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _17878_/CLK _17030_/D vssd1 vssd1 vccd1 vccd1 _17030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _14511_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ _12036_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10405_ hold4194/X _10619_/B _10404_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11385_ _12153_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__or2_1
X_14173_ hold1043/X _14198_/B _14172_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _14173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ hold3636/X _13123_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__mux2_1
X_10336_ hold4285/X _10640_/B _10335_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _17523_/Q _13056_/C _13055_/C _17522_/Q vssd1 vssd1 vccd1 vccd1 _13308_/S
+ sky130_fd_sc_hd__or4b_4
X_10267_ hold3247/X _10649_/B _10266_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10267_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _18033_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
X_12006_ _12210_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__or2_1
X_17863_ _17895_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ hold4143/X _10580_/B _10197_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10198_/X
+ sky130_fd_sc_hd__o211a_1
X_16814_ _18337_/CLK _16814_/D vssd1 vssd1 vccd1 vccd1 _16814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17794_ _17827_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ _18461_/CLK _16745_/D vssd1 vssd1 vccd1 vccd1 _16745_/Q sky130_fd_sc_hd__dfxtp_1
X_13957_ hold1561/X _13980_/B _13956_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _13957_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_199_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18063_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12908_ hold3001/X _12907_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12908_/X sky130_fd_sc_hd__mux2_1
X_16676_ _18204_/CLK _16676_/D vssd1 vssd1 vccd1 vccd1 _16676_/Q sky130_fd_sc_hd__dfxtp_1
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18415_ _18415_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_15627_ _17128_/CLK _15627_/D vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12839_ hold3065/X _12838_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12839_/X sky130_fd_sc_hd__mux2_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _18378_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ hold2695/X _15560_/A2 _15557_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _15558_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14509_ _15189_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__or2_1
X_18277_ _18334_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15489_ _15489_/A _15489_/B _15489_/C _15489_/D vssd1 vssd1 vccd1 vccd1 _15489_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08030_ hold2064/X _08029_/B _08029_/Y _08137_/A vssd1 vssd1 vccd1 vccd1 _08030_/X
+ sky130_fd_sc_hd__o211a_1
X_17228_ _17260_/CLK _17228_/D vssd1 vssd1 vccd1 vccd1 _17228_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 input30/A vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput41 input41/A vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 input60/X vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17159_ _18445_/CLK _17159_/D vssd1 vssd1 vccd1 vccd1 _17159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold825 hold859/X vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold836 hold836/A vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 hold847/A vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 input64/A sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold869 hold869/A vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08932_ hold291/X hold394/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2204 _14653_/X vssd1 vssd1 vccd1 vccd1 _18119_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2215 _12680_/X vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2226 _18199_/Q vssd1 vssd1 vccd1 vccd1 hold2226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 _14101_/X vssd1 vssd1 vccd1 vccd1 _17855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ _12426_/A _08863_/B vssd1 vssd1 vccd1 vccd1 _16050_/D sky130_fd_sc_hd__and2_1
Xhold1503 _15802_/Q vssd1 vssd1 vccd1 vccd1 hold1503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2248 _18125_/Q vssd1 vssd1 vccd1 vccd1 hold2248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 _15112_/X vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 _08444_/X vssd1 vssd1 vccd1 vccd1 _15852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 _18378_/Q vssd1 vssd1 vccd1 vccd1 hold1525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1536 _13026_/X vssd1 vssd1 vccd1 vccd1 _13028_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07814_ _15105_/A _15103_/A _15535_/A _15099_/A vssd1 vssd1 vccd1 vccd1 _07817_/B
+ sky130_fd_sc_hd__or4_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1547 _14404_/X vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08794_ _15482_/A hold292/X vssd1 vssd1 vccd1 vccd1 _16017_/D sky130_fd_sc_hd__and2_1
Xhold1558 _14739_/X vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1569 _18026_/Q vssd1 vssd1 vccd1 vccd1 hold1569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09415_ _07804_/A _09456_/B _15334_/A _09414_/X vssd1 vssd1 vccd1 vccd1 _09415_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09346_ hold173/A hold335/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__or3_1
XFILLER_0_48_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _15553_/A hold2290/X _09277_/S vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ _08504_/A hold607/X vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__and2_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ _12301_/A _11170_/B vssd1 vssd1 vccd1 vccd1 _11170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4140 _13351_/X vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10121_ hold1887/X hold3179/X _10481_/S vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__mux2_1
Xhold4151 _16643_/Q vssd1 vssd1 vccd1 vccd1 hold4151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4162 _13414_/X vssd1 vssd1 vccd1 vccd1 _17591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4173 _11908_/X vssd1 vssd1 vccd1 vccd1 _17126_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4184 _17221_/Q vssd1 vssd1 vccd1 vccd1 hold4184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4195 _10405_/X vssd1 vssd1 vccd1 vccd1 _16625_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3450 _17437_/Q vssd1 vssd1 vccd1 vccd1 hold3450/X sky130_fd_sc_hd__dlygate4sd3_1
X_10052_ _16508_/Q _10070_/B _10271_/S vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__and3_1
Xhold3461 _17262_/Q vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3472 _17428_/Q vssd1 vssd1 vccd1 vccd1 hold3472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3483 _13753_/X vssd1 vssd1 vccd1 vccd1 _17704_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3494 _12806_/X vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2760 _17998_/Q vssd1 vssd1 vccd1 vccd1 hold2760/X sky130_fd_sc_hd__dlygate4sd3_1
X_14860_ _14984_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__or2_1
Xhold2771 _18304_/Q vssd1 vssd1 vccd1 vccd1 hold2771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2782 _08451_/X vssd1 vssd1 vccd1 vccd1 _15854_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2793 _18159_/Q vssd1 vssd1 vccd1 vccd1 hold2793/X sky130_fd_sc_hd__dlygate4sd3_1
X_13811_ _17724_/Q _13811_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _13811_/X sky130_fd_sc_hd__and3_1
XFILLER_0_187_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14791_ hold2274/X _14822_/B _14790_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14791_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_292_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16530_ _18126_/CLK _16530_/D vssd1 vssd1 vccd1 vccd1 _16530_/Q sky130_fd_sc_hd__dfxtp_1
X_13742_ hold2854/X hold4526/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13743_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10954_ hold4451/X _11726_/B _10953_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_221_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17904_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16461_ _18420_/CLK _16461_/D vssd1 vssd1 vccd1 vccd1 _16461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ hold2637/X hold3344/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13674_/B sky130_fd_sc_hd__mux2_1
X_10885_ hold4234/X _11171_/B _10884_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10885_/X
+ sky130_fd_sc_hd__o211a_1
X_18200_ _18218_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _15489_/A _15412_/B _15412_/C _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_94_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12624_ _12855_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _17384_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16392_ _18273_/CLK _16392_/D vssd1 vssd1 vccd1 vccd1 _16392_/Q sky130_fd_sc_hd__dfxtp_1
X_18131_ _18131_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15343_ _15490_/A1 _15335_/X _15342_/X _15490_/B1 hold5825/A vssd1 vssd1 vccd1 vccd1
+ _15343_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12555_ _12924_/A _12555_/B vssd1 vssd1 vccd1 vccd1 _17361_/D sky130_fd_sc_hd__and2_1
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ hold4277/X _11792_/B _11505_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__o211a_1
X_18062_ _18062_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
X_15274_ _15374_/A _15274_/B vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ _17336_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ _17893_/CLK _17013_/D vssd1 vssd1 vccd1 vccd1 _17013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14225_ hold5968/X _14216_/Y hold668/X _14368_/A vssd1 vssd1 vccd1 vccd1 hold669/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ hold4367/X _11726_/B _11436_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ hold799/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14156_/X sky130_fd_sc_hd__or2_1
X_11368_ hold5435/X _11753_/B _11367_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11368_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13106_/X _16906_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
X_10319_ hold1836/X _16597_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__mux2_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ hold1322/X _14094_/B _14086_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14087_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ hold4585/X _12323_/B _11298_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13048_/A _13034_/X _13046_/A vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__a21o_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _18043_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _17877_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_309_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14989_ hold2272/X _15004_/B _14988_/X _15364_/A vssd1 vssd1 vccd1 vccd1 _14989_/X
+ sky130_fd_sc_hd__o211a_1
X_17777_ _17777_/CLK _17777_/D vssd1 vssd1 vccd1 vccd1 _17777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ _18222_/CLK _16728_/D vssd1 vssd1 vccd1 vccd1 _16728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16659_ _18185_/CLK _16659_/D vssd1 vssd1 vccd1 vccd1 _16659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09200_ _15529_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09131_ hold2953/X _09177_/A2 _09130_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09131_/X
+ sky130_fd_sc_hd__o211a_1
X_18329_ _18330_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ hold291/X hold397/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _15527_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08013_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold600 hold600/A vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 hold611/A vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold622 hold622/A vssd1 vssd1 vccd1 vccd1 input55/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold633/A vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold644 hold644/A vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 hold655/A vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__clkbuf_4
Xhold666 input62/X vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__buf_1
Xhold677 hold677/A vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/A vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 hold699/A vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ hold5619/X _10780_/A2 _09963_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _09964_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2001 _15108_/X vssd1 vssd1 vccd1 vccd1 _18338_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 _18065_/Q vssd1 vssd1 vccd1 vccd1 hold2012/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08915_ _12426_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _16075_/D sky130_fd_sc_hd__and2_1
Xhold2023 _14823_/X vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09895_ _09989_/A _09998_/B _09894_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09895_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2034 _15845_/Q vssd1 vssd1 vccd1 vccd1 hold2034/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _07973_/X vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1300 _17997_/Q vssd1 vssd1 vccd1 vccd1 hold1300/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _16275_/Q vssd1 vssd1 vccd1 vccd1 hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2056 _18158_/Q vssd1 vssd1 vccd1 vccd1 hold2056/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 _17848_/Q vssd1 vssd1 vccd1 vccd1 hold1322/X sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ hold8/X hold190/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__mux2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2067 _14095_/X vssd1 vssd1 vccd1 vccd1 _17852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1333 _15124_/X vssd1 vssd1 vccd1 vccd1 _18346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 _18368_/Q vssd1 vssd1 vccd1 vccd1 hold2078/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 _18163_/Q vssd1 vssd1 vccd1 vccd1 hold1344/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2089 _08501_/X vssd1 vssd1 vccd1 vccd1 _15879_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1355 _16217_/Q vssd1 vssd1 vccd1 vccd1 hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1366 _15832_/Q vssd1 vssd1 vccd1 vccd1 hold1366/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1377 _17793_/Q vssd1 vssd1 vccd1 vccd1 hold1377/X sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ hold149/X _16009_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__mux2_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1388 _08288_/X vssd1 vssd1 vccd1 vccd1 _15777_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _18023_/Q vssd1 vssd1 vccd1 vccd1 hold1399/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ hold1872/X hold3616/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _15551_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _12343_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ hold4530/X _13844_/B _12270_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _12271_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14010_ _14511_/A _14050_/B vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__or2_1
X_11222_ _16898_/Q _11222_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__and3_1
X_11153_ _16875_/Q _11156_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__and3_1
X_10104_ _10527_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__or2_1
X_15961_ _16128_/CLK _15961_/D vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__dfxtp_1
X_11084_ hold1424/X _16852_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__mux2_1
Xhold3280 _10669_/X vssd1 vssd1 vccd1 vccd1 _16713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3291 _17686_/Q vssd1 vssd1 vccd1 vccd1 hold3291/X sky130_fd_sc_hd__dlygate4sd3_1
X_17700_ _17732_/CLK _17700_/D vssd1 vssd1 vccd1 vccd1 _17700_/Q sky130_fd_sc_hd__dfxtp_1
X_14912_ _14913_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__nor2_2
X_10035_ _13206_/A _10380_/A _10034_/X vssd1 vssd1 vccd1 vccd1 _10035_/Y sky130_fd_sc_hd__a21oi_1
X_15892_ _17314_/CLK _15892_/D vssd1 vssd1 vccd1 vccd1 hold640/A sky130_fd_sc_hd__dfxtp_1
Xhold2590 _16199_/Q vssd1 vssd1 vccd1 vccd1 hold2590/X sky130_fd_sc_hd__dlygate4sd3_1
X_17631_ _17697_/CLK _17631_/D vssd1 vssd1 vccd1 vccd1 _17631_/Q sky130_fd_sc_hd__dfxtp_1
X_14843_ _14843_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14864_/B sky130_fd_sc_hd__or2_4
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ _17722_/CLK _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14774_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__nand2_1
X_11986_ hold3347/X _12374_/B _11985_/X _12274_/C1 vssd1 vssd1 vccd1 vccd1 _11986_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16513_ _18330_/CLK _16513_/D vssd1 vssd1 vccd1 vccd1 _16513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13725_ _13734_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__or2_1
X_10937_ hold2324/X hold4248/X _11765_/C vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__mux2_1
X_17493_ _17506_/CLK _17493_/D vssd1 vssd1 vccd1 vccd1 _17493_/Q sky130_fd_sc_hd__dfxtp_1
X_16444_ _18389_/CLK _16444_/D vssd1 vssd1 vccd1 vccd1 _16444_/Q sky130_fd_sc_hd__dfxtp_1
X_13656_ _13758_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ hold1722/X _16780_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ hold2656/X _17380_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__mux2_1
X_16375_ _18390_/CLK _16375_/D vssd1 vssd1 vccd1 vccd1 _16375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13788_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ hold1002/X _16757_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__mux2_1
X_18114_ _18210_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
X_15326_ _17336_/Q _09362_/C _15485_/B1 hold361/X vssd1 vssd1 vccd1 vccd1 _15326_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12538_ hold1471/X hold3581/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18045_ _18047_/CLK _18045_/D vssd1 vssd1 vccd1 vccd1 _18045_/Q sky130_fd_sc_hd__dfxtp_1
X_15257_ _16134_/Q _09357_/A _15484_/B1 hold293/X _15256_/X vssd1 vssd1 vccd1 vccd1
+ _15262_/B sky130_fd_sc_hd__a221o_1
X_12469_ hold2/X _08598_/B _08999_/B _12468_/X _15414_/A vssd1 vssd1 vccd1 vccd1 hold3/A
+ sky130_fd_sc_hd__o311a_1
Xhold4909 _17264_/Q vssd1 vssd1 vccd1 vccd1 hold4909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14208_ _14726_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__or2_1
X_15188_ hold5958/X _15219_/B _15187_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14139_ hold829/X hold587/X _14138_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 hold830/A
+ sky130_fd_sc_hd__o211a_1
Xfanout409 _14280_/B vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__clkbuf_8
X_08700_ _15344_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _15971_/D sky130_fd_sc_hd__and2_1
X_09680_ hold1614/X _16384_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_143_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18266_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08631_ hold214/X hold409/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08632_/B sky130_fd_sc_hd__mux2_1
X_17829_ _17829_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ hold179/X hold181/X _08562_/S vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__mux2_1
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ hold1240/X _08486_/B _08492_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08493_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ hold800/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09045_ _12442_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _16139_/D sky130_fd_sc_hd__and2_1
XFILLER_0_128_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold441/A vssd1 vssd1 vccd1 vccd1 input36/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 hold452/A vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 la_data_in[15] vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 hold485/A vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold496 hold496/A vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 hold799/X vssd1 vssd1 vccd1 vccd1 _14728_/A sky130_fd_sc_hd__buf_8
Xfanout921 hold730/X vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__clkbuf_16
X_09947_ hold1401/X _16473_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__mux2_1
Xfanout932 hold734/X vssd1 vssd1 vccd1 vccd1 hold735/A sky130_fd_sc_hd__buf_6
Xfanout943 hold747/X vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__clkbuf_16
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ hold1391/X hold4291/X _10271_/S vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__mux2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _16187_/Q vssd1 vssd1 vccd1 vccd1 hold1130/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _09071_/X vssd1 vssd1 vccd1 vccd1 _16150_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _12438_/A hold504/X vssd1 vssd1 vccd1 vccd1 _16033_/D sky130_fd_sc_hd__and2_1
Xhold1152 _18204_/Q vssd1 vssd1 vccd1 vccd1 hold1152/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _15640_/Q vssd1 vssd1 vccd1 vccd1 hold1163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 _15721_/Q vssd1 vssd1 vccd1 vccd1 hold1174/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _16191_/Q vssd1 vssd1 vccd1 vccd1 hold1185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _14464_/X vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ hold2354/X hold3805/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _17081_/Q _12338_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13510_ hold4117/X _13814_/B _13509_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _11106_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__or2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ hold2246/X _14487_/B _14489_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _14490_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ hold3357/X _13823_/B _13440_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _17600_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _11076_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _17981_/CLK _16160_/D vssd1 vssd1 vccd1 vccd1 _16160_/Q sky130_fd_sc_hd__dfxtp_1
X_13372_ hold5122/X _13886_/B _13371_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13372_/X
+ sky130_fd_sc_hd__o211a_1
X_10584_ hold3852/X _10491_/A _10583_/X vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__a21oi_1
X_15111_ _15219_/A _15113_/B vssd1 vssd1 vccd1 vccd1 _15111_/Y sky130_fd_sc_hd__nand2_1
X_12323_ _17265_/Q _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and3_1
X_16091_ _18406_/CLK _16091_/D vssd1 vssd1 vccd1 vccd1 hold598/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15042_ _15394_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12254_ hold1736/X hold5019/X _13388_/S vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__mux2_1
X_11205_ hold5260/X _11658_/A _11204_/X vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12185_ hold2010/X hold4486/X _12377_/C vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__mux2_1
X_11136_ _11136_/A _11136_/B vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__or2_1
X_16993_ _17873_/CLK _16993_/D vssd1 vssd1 vccd1 vccd1 _16993_/Q sky130_fd_sc_hd__dfxtp_1
X_15944_ _18406_/CLK _15944_/D vssd1 vssd1 vccd1 vccd1 hold712/A sky130_fd_sc_hd__dfxtp_1
X_11067_ _11067_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__or2_1
X_10018_ _11155_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10018_/Y sky130_fd_sc_hd__nor2_1
X_15875_ _17747_/CLK _15875_/D vssd1 vssd1 vccd1 vccd1 _15875_/Q sky130_fd_sc_hd__dfxtp_1
X_14826_ _15219_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14826_/Y sky130_fd_sc_hd__nand2_1
X_17614_ _17678_/CLK _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _18360_/CLK _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_1
X_14757_ hold2300/X _14772_/B _14756_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14757_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ hold2326/X hold3521/X _12356_/C vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ hold4811/X _13805_/B _13707_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13708_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17476_ _17785_/CLK _17476_/D vssd1 vssd1 vccd1 vccd1 _17476_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _15189_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16427_ _18380_/CLK _16427_/D vssd1 vssd1 vccd1 vccd1 _16427_/Q sky130_fd_sc_hd__dfxtp_1
X_13639_ hold4283/X _13814_/B _13638_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _17666_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16358_ _18337_/CLK _16358_/D vssd1 vssd1 vccd1 vccd1 _16358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ hold723/X _09365_/B _09392_/C hold648/X _15308_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5407 _16799_/Q vssd1 vssd1 vccd1 vccd1 hold5407/X sky130_fd_sc_hd__dlygate4sd3_1
X_16289_ _18409_/CLK _16289_/D vssd1 vssd1 vccd1 vccd1 _16289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5418 _10792_/X vssd1 vssd1 vccd1 vccd1 _16754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5429 _16493_/Q vssd1 vssd1 vccd1 vccd1 hold5429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4706 _16592_/Q vssd1 vssd1 vccd1 vccd1 hold4706/X sky130_fd_sc_hd__dlygate4sd3_1
X_18028_ _18208_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4717 _10813_/X vssd1 vssd1 vccd1 vccd1 _16761_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4728 _11842_/X vssd1 vssd1 vccd1 vccd1 _17104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4739 _17192_/Q vssd1 vssd1 vccd1 vccd1 hold4739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout206 _11222_/B vssd1 vssd1 vccd1 vccd1 _11789_/B sky130_fd_sc_hd__buf_4
Xfanout217 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__clkbuf_4
X_09801_ _10779_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__or2_1
Xfanout228 _10897_/A2 vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__buf_4
XFILLER_0_157_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout239 _10601_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__clkbuf_8
X_07993_ _08504_/A _14681_/A vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_2
X_09732_ _09924_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09663_ _09975_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08614_ _09021_/A _08614_/B vssd1 vssd1 vccd1 vccd1 _15929_/D sky130_fd_sc_hd__and2_1
X_09594_ _10506_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08545_ _12442_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _15896_/D sky130_fd_sc_hd__and2_1
XFILLER_0_166_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _14529_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5930 _17555_/Q vssd1 vssd1 vccd1 vccd1 hold5930/X sky130_fd_sc_hd__dlygate4sd3_1
X_09028_ hold71/X hold670/X _09028_/S vssd1 vssd1 vccd1 vccd1 hold671/A sky130_fd_sc_hd__mux2_1
Xhold5941 hold6004/X vssd1 vssd1 vccd1 vccd1 hold5941/X sky130_fd_sc_hd__buf_1
XFILLER_0_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5952 _18241_/Q vssd1 vssd1 vccd1 vccd1 hold5952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5963 _18007_/Q vssd1 vssd1 vccd1 vccd1 hold5963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5974 _15848_/Q vssd1 vssd1 vccd1 vccd1 hold5974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5985 data_in[20] vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5996 _18404_/Q vssd1 vssd1 vccd1 vccd1 hold5996/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__buf_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__buf_4
Xfanout751 _13909_/A vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__buf_4
Xfanout762 fanout763/X vssd1 vssd1 vccd1 vccd1 _14402_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout773 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _13792_/C1 sky130_fd_sc_hd__buf_4
X_13990_ _14330_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13990_/X sky130_fd_sc_hd__or2_1
Xfanout784 _14203_/C1 vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__buf_4
Xfanout795 _15060_/A vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__buf_4
XFILLER_0_172_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ hold3593/X _12940_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12942_/B sky130_fd_sc_hd__mux2_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _17583_/CLK _15660_/D vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ hold3281/X _12871_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__mux2_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _14850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ hold2405/X _14610_/B _14610_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14611_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _12210_/A _11823_/B vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__or2_1
XANTENNA_133 hold5983/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _17216_/CLK _15591_/D vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _18410_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _17330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ hold2312/X _14541_/B _14541_/Y _14390_/A vssd1 vssd1 vccd1 vccd1 _14542_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ hold5233/X _11658_/A _11753_/X vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17718_/CLK _17261_/D vssd1 vssd1 vccd1 vccd1 _17261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ hold5462/X _11216_/B _10704_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14473_ _15099_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14473_/X sky130_fd_sc_hd__or2_1
X_11685_ _12036_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__or2_1
X_16212_ _17435_/CLK _16212_/D vssd1 vssd1 vccd1 vccd1 _16212_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ hold1366/X hold3396/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13425_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ _17692_/CLK _17192_/D vssd1 vssd1 vccd1 vccd1 _17192_/Q sky130_fd_sc_hd__dfxtp_1
X_10636_ _11218_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16143_ _17314_/CLK _16143_/D vssd1 vssd1 vccd1 vccd1 hold477/A sky130_fd_sc_hd__dfxtp_1
X_13355_ hold1128/X hold3894/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__mux2_1
X_10567_ _11194_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ hold3950/X _12018_/A _12305_/X vssd1 vssd1 vccd1 vccd1 _12306_/Y sky130_fd_sc_hd__a21oi_1
X_16074_ _18421_/CLK _16074_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13286_ _13286_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10498_ _10592_/A _10646_/B _10497_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _16656_/D
+ sky130_fd_sc_hd__o211a_1
X_15025_ _15187_/A hold1348/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15026_/B sky130_fd_sc_hd__mux2_1
X_12237_ _12255_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12168_ _12255_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11119_ hold5474/X _11213_/B _11118_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12099_ _13797_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
X_16976_ _17856_/CLK _16976_/D vssd1 vssd1 vccd1 vccd1 _16976_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 input6/A vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _17530_/CLK _15927_/D vssd1 vssd1 vccd1 vccd1 hold551/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _17741_/CLK _15858_/D vssd1 vssd1 vccd1 vccd1 _15858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ hold1292/X _14822_/B _14808_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14809_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789_ _17725_/CLK _15789_/D vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08330_ hold2199/X _08336_/A2 _08329_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08330_/X
+ sky130_fd_sc_hd__o211a_1
X_17528_ _17528_/CLK _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ hold1501/X _08262_/B _08260_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08261_/X
+ sky130_fd_sc_hd__o211a_1
X_17459_ _18458_/CLK _17459_/D vssd1 vssd1 vccd1 vccd1 _17459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08192_ hold1414/X _08213_/B _08191_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _08192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5204 _13501_/X vssd1 vssd1 vccd1 vccd1 _17620_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5215 _17740_/Q vssd1 vssd1 vccd1 vccd1 hold5215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5226 _10012_/Y vssd1 vssd1 vccd1 vccd1 _16494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5237 _11772_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4503 _12136_/X vssd1 vssd1 vccd1 vccd1 _17202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5248 _16736_/Q vssd1 vssd1 vccd1 vccd1 hold5248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5259 _10006_/Y vssd1 vssd1 vccd1 vccd1 _16492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4514 _16984_/Q vssd1 vssd1 vccd1 vccd1 hold4514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4525 _11263_/X vssd1 vssd1 vccd1 vccd1 _16911_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4536 _17249_/Q vssd1 vssd1 vccd1 vccd1 hold4536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3802 _16354_/Q vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4547 _16744_/Q vssd1 vssd1 vccd1 vccd1 hold4547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4558 _13525_/X vssd1 vssd1 vccd1 vccd1 _17628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3813 _12301_/Y vssd1 vssd1 vccd1 vccd1 _17257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3824 _13870_/Y vssd1 vssd1 vccd1 vccd1 _17743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4569 _17137_/Q vssd1 vssd1 vccd1 vccd1 hold4569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3835 _17105_/Q vssd1 vssd1 vccd1 vccd1 hold3835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3846 _17573_/Q vssd1 vssd1 vccd1 vccd1 hold3846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3857 _16491_/Q vssd1 vssd1 vccd1 vccd1 hold3857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3868 _17113_/Q vssd1 vssd1 vccd1 vccd1 hold3868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3879 _12343_/Y vssd1 vssd1 vccd1 vccd1 _17271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07976_ _15545_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07976_/Y sky130_fd_sc_hd__nand2_1
X_09715_ hold3863/X _10001_/B _09714_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__o211a_1
X_09646_ hold3378/X _09952_/A2 _09645_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _09646_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ hold5100/X _10601_/B _09576_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ hold407/X hold513/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08459_ hold1210/X _08488_/B _08458_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08459_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ hold5403/X _11762_/B _11469_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _11470_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ hold1330/X _16631_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_246_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13140_ hold5312/X _13139_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__mux2_1
X_10352_ hold1403/X hold4365/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5760 output82/X vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_12
X_13071_ _13183_/A1 _13069_/X _13070_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13071_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_104_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5771 hold5914/X vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10283_ hold2832/X _16585_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__mux2_1
Xhold5782 output88/X vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_12
Xhold5793 hold5924/X vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__dlygate4sd3_1
X_12022_ hold4696/X _12308_/B _12021_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12022_/X
+ sky130_fd_sc_hd__o211a_1
X_16830_ _18065_/CLK _16830_/D vssd1 vssd1 vccd1 vccd1 _16830_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout570 _07991_/A2 vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__clkbuf_8
Xfanout581 hold655/X vssd1 vssd1 vccd1 vccd1 hold656/A sky130_fd_sc_hd__clkbuf_2
Xfanout592 _12814_/S vssd1 vssd1 vccd1 vccd1 _12820_/S sky130_fd_sc_hd__buf_6
X_13973_ hold1377/X _13980_/B _13972_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _13973_/X
+ sky130_fd_sc_hd__o211a_1
X_16761_ _18055_/CLK _16761_/D vssd1 vssd1 vccd1 vccd1 _16761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15712_ _17279_/CLK _15712_/D vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfxtp_1
X_12924_ _12924_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _17484_/D sky130_fd_sc_hd__and2_1
X_16692_ _18218_/CLK _16692_/D vssd1 vssd1 vccd1 vccd1 _16692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18431_ _18431_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
X_15643_ _17281_/CLK _15643_/D vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfxtp_1
X_12855_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _17461_/D sky130_fd_sc_hd__and2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ hold5158/X _12305_/B _11805_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11806_/X
+ sky130_fd_sc_hd__o211a_1
X_18362_ _18396_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ _17274_/CLK _15574_/D vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12786_ _12789_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _17438_/D sky130_fd_sc_hd__and2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17313_ _17313_/CLK _17313_/D vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _15205_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _12301_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18293_ _18315_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17244_ _17276_/CLK _17244_/D vssd1 vssd1 vccd1 vccd1 _17244_/Q sky130_fd_sc_hd__dfxtp_1
X_14456_ hold2903/X _14481_/B _14455_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _14456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ hold5689/X _11762_/B _11667_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11668_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ _13791_/A _13407_/B vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ _10619_/A _10619_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__and3_1
X_17175_ _17779_/CLK _17175_/D vssd1 vssd1 vccd1 vccd1 _17175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14387_ _14728_/A hold2287/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14388_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ hold5743/X _11789_/B _11598_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11599_/X
+ sky130_fd_sc_hd__o211a_1
X_16126_ _17342_/CLK _16126_/D vssd1 vssd1 vccd1 vccd1 hold714/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13338_ _13767_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16057_ _17331_/CLK _16057_/D vssd1 vssd1 vccd1 vccd1 _16057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13269_ _13268_/X hold3630/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__mux2_1
Xhold3109 _17468_/Q vssd1 vssd1 vccd1 vccd1 hold3109/X sky130_fd_sc_hd__dlygate4sd3_1
X_15008_ hold730/X _15012_/B vssd1 vssd1 vccd1 vccd1 _15008_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2408 _15534_/X vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2419 _18177_/Q vssd1 vssd1 vccd1 vccd1 hold2419/X sky130_fd_sc_hd__dlygate4sd3_1
X_07830_ _14843_/A hold816/X vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__or2_4
Xhold1707 _14797_/X vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1718 _18395_/Q vssd1 vssd1 vccd1 vccd1 hold1718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 hold5832/X vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__clkbuf_4
X_16959_ _17829_/CLK _16959_/D vssd1 vssd1 vccd1 vccd1 _16959_/Q sky130_fd_sc_hd__dfxtp_1
X_09500_ hold1932/X _13062_/A _09998_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _07785_/Y hold681/X _15314_/A _09430_/X vssd1 vssd1 vccd1 vccd1 hold682/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _09362_/A _09392_/B _09362_/C _09362_/D vssd1 vssd1 vccd1 vccd1 _09369_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _15537_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08313_/X sky130_fd_sc_hd__or2_1
XFILLER_0_176_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09293_ _15515_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__or2_1
XANTENNA_11 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _14517_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08244_/X sky130_fd_sc_hd__or2_1
XANTENNA_33 fanout337/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_44 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 _15535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 hold335/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_77 hold883/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _14218_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__or2_1
XANTENNA_88 hold5830/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_99 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5001 _17252_/Q vssd1 vssd1 vccd1 vccd1 hold5001/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5012 _10123_/X vssd1 vssd1 vccd1 vccd1 _16531_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5023 _17211_/Q vssd1 vssd1 vccd1 vccd1 hold5023/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5034 _17229_/Q vssd1 vssd1 vccd1 vccd1 hold5034/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4300 _10414_/X vssd1 vssd1 vccd1 vccd1 _16628_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5045 _12169_/X vssd1 vssd1 vccd1 vccd1 _17213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4311 _17126_/Q vssd1 vssd1 vccd1 vccd1 hold4311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5056 _16376_/Q vssd1 vssd1 vccd1 vccd1 hold5056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4322 _10222_/X vssd1 vssd1 vccd1 vccd1 _16564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5067 _13465_/X vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput140 hold5820/X vssd1 vssd1 vccd1 vccd1 hold5821/A sky130_fd_sc_hd__buf_6
Xhold4333 _17690_/Q vssd1 vssd1 vccd1 vccd1 hold4333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5078 _17244_/Q vssd1 vssd1 vccd1 vccd1 hold5078/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4344 _12016_/X vssd1 vssd1 vccd1 vccd1 _17162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5089 _11923_/X vssd1 vssd1 vccd1 vccd1 _17131_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4355 _17065_/Q vssd1 vssd1 vccd1 vccd1 hold4355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3610 _16711_/Q vssd1 vssd1 vccd1 vccd1 hold3610/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_101_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3621 _10618_/Y vssd1 vssd1 vccd1 vccd1 _16696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4366 _10258_/X vssd1 vssd1 vccd1 vccd1 _16576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4377 _17613_/Q vssd1 vssd1 vccd1 vccd1 hold4377/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3632 _10636_/Y vssd1 vssd1 vccd1 vccd1 _16702_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4388 _10513_/X vssd1 vssd1 vccd1 vccd1 _16661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3643 _10644_/Y vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4399 _17057_/Q vssd1 vssd1 vccd1 vccd1 hold4399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3654 _16342_/Q vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3665 _16717_/Q vssd1 vssd1 vccd1 vccd1 hold3665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2920 _17973_/Q vssd1 vssd1 vccd1 vccd1 hold2920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2931 _14699_/X vssd1 vssd1 vccd1 vccd1 _18141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3676 _10059_/Y vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2942 _18299_/Q vssd1 vssd1 vccd1 vccd1 hold2942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3687 _17567_/Q vssd1 vssd1 vccd1 vccd1 hold3687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2953 _16178_/Q vssd1 vssd1 vccd1 vccd1 hold2953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3698 _11170_/Y vssd1 vssd1 vccd1 vccd1 _16880_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 _07945_/X vssd1 vssd1 vccd1 vccd1 _15615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2975 _17835_/Q vssd1 vssd1 vccd1 vccd1 hold2975/X sky130_fd_sc_hd__dlygate4sd3_1
X_07959_ hold2789/X _07991_/A2 _07958_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07959_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2986 _14460_/X vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2997 _15778_/Q vssd1 vssd1 vccd1 vccd1 hold2997/X sky130_fd_sc_hd__dlygate4sd3_1
X_10970_ hold1154/X hold3948/X _11066_/S vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__mux2_1
X_09629_ hold2272/X _16367_/Q _09893_/S vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ hold2548/X _17391_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ hold2951/X _17368_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__mux2_1
X_14310_ _15205_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__or2_1
X_11522_ hold1686/X _16998_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__mux2_1
X_15290_ hold390/X _15486_/A2 _15446_/B1 _16058_/Q vssd1 vssd1 vccd1 vccd1 _15290_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ hold2936/X _14266_/B _14240_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _14241_/X
+ sky130_fd_sc_hd__o211a_1
X_11453_ hold1939/X hold3408/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10404_ _10524_/A _10404_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__or2_1
X_14172_ _14511_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14172_/X sky130_fd_sc_hd__or2_1
X_11384_ hold2355/X _16952_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__mux2_1
X_13123_ _13122_/X hold5893/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__mux2_1
X_10335_ _10554_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/X sky130_fd_sc_hd__or2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13197_/S
+ sky130_fd_sc_hd__and4b_4
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5590 _16709_/Q vssd1 vssd1 vccd1 vccd1 hold5590/X sky130_fd_sc_hd__dlygate4sd3_1
X_17931_ _18228_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
X_10266_ _10554_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ hold2471/X hold3230/X _12308_/C vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17862_ _17862_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10197_ _10548_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16813_ _18305_/CLK _16813_/D vssd1 vssd1 vccd1 vccd1 _16813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17793_ _17889_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_1
X_16744_ _18043_/CLK _16744_/D vssd1 vssd1 vccd1 vccd1 _16744_/Q sky130_fd_sc_hd__dfxtp_1
X_13956_ _15517_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ hold1917/X _17480_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__mux2_1
X_16675_ _18233_/CLK _16675_/D vssd1 vssd1 vccd1 vccd1 _16675_/Q sky130_fd_sc_hd__dfxtp_1
X_13887_ hold3185/X _13779_/A _13886_/X vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ _18414_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15626_ _17592_/CLK _15626_/D vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfxtp_1
X_12838_ hold2652/X _17457_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ _18391_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_12769_ hold2536/X _17434_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15557_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18216_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14508_ hold2705/X _14554_/A2 _14507_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _14508_/X
+ sky130_fd_sc_hd__o211a_1
X_15488_ hold704/X _09392_/C _15485_/X vssd1 vssd1 vccd1 vccd1 _15489_/D sky130_fd_sc_hd__a21o_1
X_18276_ _18308_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 input20/A vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17227_ _17227_/CLK _17227_/D vssd1 vssd1 vccd1 vccd1 _17227_/Q sky130_fd_sc_hd__dfxtp_1
Xinput31 input31/A vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14439_ hold770/X _14445_/B vssd1 vssd1 vccd1 vccd1 hold771/A sky130_fd_sc_hd__or2_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 input42/A vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 input53/A vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 input64/A vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
X_17158_ _17592_/CLK _17158_/D vssd1 vssd1 vccd1 vccd1 _17158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 hold815/A vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__buf_6
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold837 hold837/A vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _17522_/CLK _16109_/D vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__dfxtp_1
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ hold2346/X _16484_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__mux2_1
X_17089_ _17777_/CLK _17089_/D vssd1 vssd1 vccd1 vccd1 _17089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold859 input64/X vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ _12442_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _16083_/D sky130_fd_sc_hd__and2_1
XFILLER_0_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2205 _16227_/Q vssd1 vssd1 vccd1 vccd1 hold2205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2216 _15743_/Q vssd1 vssd1 vccd1 vccd1 hold2216/X sky130_fd_sc_hd__dlygate4sd3_1
X_08862_ hold380/X hold400/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08863_/B sky130_fd_sc_hd__mux2_1
Xhold2227 _14819_/X vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2238 _16233_/Q vssd1 vssd1 vccd1 vccd1 hold2238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _14665_/X vssd1 vssd1 vccd1 vccd1 _18125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 _16287_/Q vssd1 vssd1 vccd1 vccd1 hold1504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1515 _18134_/Q vssd1 vssd1 vccd1 vccd1 hold1515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _15192_/X vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ _15531_/A _14988_/A _14986_/A _14984_/A vssd1 vssd1 vccd1 vccd1 _07817_/A
+ sky130_fd_sc_hd__or4_1
Xhold1537 _13028_/X vssd1 vssd1 vccd1 vccd1 _17519_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08793_ hold291/X _16017_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__mux2_1
Xhold1548 _15634_/Q vssd1 vssd1 vccd1 vccd1 hold1548/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1559 _18224_/Q vssd1 vssd1 vccd1 vccd1 hold1559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09414_ _09438_/B _16293_/Q vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ hold800/X hold770/X _15551_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09359_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_30_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _12756_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _16249_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ hold279/X hold606/A hold298/A hold624/A vssd1 vssd1 vccd1 vccd1 hold607/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_105_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _14218_/A hold2396/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08089_ hold2469/X _08088_/B _08088_/Y _13941_/A vssd1 vssd1 vccd1 vccd1 _08089_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4130 _10249_/X vssd1 vssd1 vccd1 vccd1 _16573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4141 _16621_/Q vssd1 vssd1 vccd1 vccd1 hold4141/X sky130_fd_sc_hd__dlygate4sd3_1
X_10120_ hold4246/X _10643_/B _10119_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10120_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4152 _10363_/X vssd1 vssd1 vccd1 vccd1 _16611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4163 _17631_/Q vssd1 vssd1 vccd1 vccd1 hold4163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4174 _16704_/Q vssd1 vssd1 vccd1 vccd1 hold4174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3440 _17020_/Q vssd1 vssd1 vccd1 vccd1 hold3440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4185 _12097_/X vssd1 vssd1 vccd1 vccd1 _17189_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10051_ _10588_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _16507_/D sky130_fd_sc_hd__nor2_1
Xhold4196 _16653_/Q vssd1 vssd1 vccd1 vccd1 hold4196/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3451 _17508_/Q vssd1 vssd1 vccd1 vccd1 hold3451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3462 _12220_/X vssd1 vssd1 vccd1 vccd1 _17230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3473 _12755_/X vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3484 _16385_/Q vssd1 vssd1 vccd1 vccd1 hold3484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2750 _16226_/Q vssd1 vssd1 vccd1 vccd1 hold2750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3495 _17170_/Q vssd1 vssd1 vccd1 vccd1 hold3495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2761 _14400_/X vssd1 vssd1 vccd1 vccd1 _17998_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2772 _15755_/Q vssd1 vssd1 vccd1 vccd1 hold2772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2783 _17891_/Q vssd1 vssd1 vccd1 vccd1 hold2783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2794 _14737_/X vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13810_ _13822_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13810_/Y sky130_fd_sc_hd__nor2_1
X_14790_ _15129_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14790_/X sky130_fd_sc_hd__or2_1
X_13741_ hold4983/X _13856_/B _13740_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _11631_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16460_ _18334_/CLK _16460_/D vssd1 vssd1 vccd1 vccd1 _16460_/Q sky130_fd_sc_hd__dfxtp_1
X_13672_ hold3273/X _13862_/B _13671_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13672_/X
+ sky130_fd_sc_hd__o211a_1
X_10884_ _11652_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15411_ _16305_/Q _15477_/A2 _15487_/B1 _16093_/Q _15410_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/D sky130_fd_sc_hd__a221o_1
X_12623_ hold3074/X _12622_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12623_/X sky130_fd_sc_hd__mux2_1
X_16391_ _18304_/CLK _16391_/D vssd1 vssd1 vccd1 vccd1 _16391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15342_ _15489_/A _15342_/B _15342_/C _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/X
+ sky130_fd_sc_hd__or4_1
X_18130_ _18206_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_261_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17742_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12554_ hold3317/X _12553_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _11697_/A _11505_/B vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15273_ _15490_/A1 _15265_/X _15272_/X _15490_/B1 hold4842/X vssd1 vssd1 vccd1 vccd1
+ _15273_/X sky130_fd_sc_hd__a32o_1
X_18061_ _18061_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ hold17/X _08598_/B _08999_/B _12484_/X _09047_/A vssd1 vssd1 vccd1 vccd1
+ hold18/A sky130_fd_sc_hd__o311a_1
XFILLER_0_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17012_ _17862_/CLK _17012_/D vssd1 vssd1 vccd1 vccd1 _17012_/Q sky130_fd_sc_hd__dfxtp_1
X_14224_ hold667/X _14230_/B vssd1 vssd1 vccd1 vccd1 hold668/A sky130_fd_sc_hd__or2_1
X_11436_ _11631_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14155_ hold2421/X _14148_/B _14154_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _14155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11367_ _11658_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ _17564_/Q _17098_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__mux2_1
X_10318_ hold4413/X _10649_/B _10317_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10318_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ _15539_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14086_/X sky130_fd_sc_hd__or2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _12036_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__or2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _15284_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _17522_/D sky130_fd_sc_hd__and2_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _18042_/CLK hold669/X vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_1
X_10249_ hold4129/X _10631_/B _10248_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10249_/X
+ sky130_fd_sc_hd__o211a_1
X_17845_ _17877_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_1
X_17776_ _17799_/CLK _17776_/D vssd1 vssd1 vccd1 vccd1 _17776_/Q sky130_fd_sc_hd__dfxtp_1
X_14988_ _14988_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ _18158_/CLK _16727_/D vssd1 vssd1 vccd1 vccd1 _16727_/Q sky130_fd_sc_hd__dfxtp_1
X_13939_ _13939_/A _13939_/B vssd1 vssd1 vccd1 vccd1 _17777_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16658_ _18216_/CLK _16658_/D vssd1 vssd1 vccd1 vccd1 _16658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15609_ _17257_/CLK _15609_/D vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16589_ _18266_/CLK _16589_/D vssd1 vssd1 vccd1 vccd1 _16589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09130_ _15513_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__or2_1
X_18328_ _18392_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ _12426_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _16147_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18259_ _18395_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08012_ hold2471/X _08029_/B _08011_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _08012_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 hold601/A vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold612 hold612/A vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold623 input55/X vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__buf_1
XFILLER_0_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold634 hold634/A vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 hold645/A vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold656 hold656/A vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__clkbuf_8
Xhold667 hold667/A vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__buf_6
Xhold678 hold678/A vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _11106_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__or2_1
Xhold689 hold689/A vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18406_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08914_ hold140/X hold688/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2002 _18391_/Q vssd1 vssd1 vccd1 vccd1 hold2002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2013 _14538_/X vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ _09918_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__or2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _15775_/Q vssd1 vssd1 vccd1 vccd1 hold2024/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2035 _08430_/X vssd1 vssd1 vccd1 vccd1 _15845_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 _17935_/Q vssd1 vssd1 vccd1 vccd1 hold2046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1301 _14398_/X vssd1 vssd1 vccd1 vccd1 _17997_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _15454_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _16041_/D sky130_fd_sc_hd__and2_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _09330_/X vssd1 vssd1 vccd1 vccd1 _16275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2057 _14733_/X vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 _14087_/X vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2068 _18038_/Q vssd1 vssd1 vccd1 vccd1 hold2068/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 _15170_/X vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _17776_/Q vssd1 vssd1 vccd1 vccd1 hold1334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 _14745_/X vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1356 _09211_/X vssd1 vssd1 vccd1 vccd1 _16217_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _15482_/A hold481/X vssd1 vssd1 vccd1 vccd1 _16008_/D sky130_fd_sc_hd__and2_1
Xhold1367 _08404_/X vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 _13973_/X vssd1 vssd1 vccd1 vccd1 _17793_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 _18282_/Q vssd1 vssd1 vccd1 vccd1 hold1389/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09328_ hold2314/X _09325_/B _09327_/X _14360_/A vssd1 vssd1 vccd1 vccd1 _09328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _15535_/A hold1575/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12270_ _13749_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ _12343_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11221_/Y sky130_fd_sc_hd__nor2_1
X_11152_ _11155_/A _11152_/B vssd1 vssd1 vccd1 vccd1 _11152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10103_ hold2691/X _16525_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__mux2_1
X_15960_ _17302_/CLK _15960_/D vssd1 vssd1 vccd1 vccd1 _15960_/Q sky130_fd_sc_hd__dfxtp_1
X_11083_ hold4176/X _11177_/B _11082_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _11083_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3270 _17481_/Q vssd1 vssd1 vccd1 vccd1 hold3270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3281 _17467_/Q vssd1 vssd1 vccd1 vccd1 hold3281/X sky130_fd_sc_hd__dlygate4sd3_1
X_14911_ hold1899/X hold657/X _14910_/X _15354_/A vssd1 vssd1 vccd1 vccd1 _14911_/X
+ sky130_fd_sc_hd__o211a_1
X_10034_ _16502_/Q _10571_/B _10571_/C vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__and3_1
Xhold3292 _13603_/X vssd1 vssd1 vccd1 vccd1 _17654_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15891_ _17329_/CLK _15891_/D vssd1 vssd1 vccd1 vccd1 hold447/A sky130_fd_sc_hd__dfxtp_1
Xhold2580 _18058_/Q vssd1 vssd1 vccd1 vccd1 hold2580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _17726_/CLK _17630_/D vssd1 vssd1 vccd1 vccd1 _17630_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2591 _09173_/X vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14842_ _14843_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14842_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1890 _13969_/X vssd1 vssd1 vccd1 vccd1 _17791_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17561_ _17721_/CLK _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
X_14773_ hold2419/X _14772_/B _14772_/Y _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14773_/X
+ sky130_fd_sc_hd__o211a_1
X_11985_ _12279_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16512_ _18265_/CLK _16512_/D vssd1 vssd1 vccd1 vccd1 _16512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ hold2654/X hold4167/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10936_ hold4301/X _11222_/B _10935_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _10936_/X
+ sky130_fd_sc_hd__o211a_1
X_17492_ _17506_/CLK _17492_/D vssd1 vssd1 vccd1 vccd1 _17492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ _18390_/CLK _16443_/D vssd1 vssd1 vccd1 vccd1 _16443_/Q sky130_fd_sc_hd__dfxtp_1
X_13655_ hold1738/X _17672_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ hold5548/X _09992_/B _10866_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10867_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12606_ _12909_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _17378_/D sky130_fd_sc_hd__and2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ hold2811/X _17649_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16374_ _18319_/CLK _16374_/D vssd1 vssd1 vccd1 vccd1 _16374_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ hold4831/X _11192_/B _10797_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _16756_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18392_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15325_ _15325_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15325_/X sky130_fd_sc_hd__or2_1
X_12537_ _12936_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _17355_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18044_ _18047_/CLK hold955/X vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__dfxtp_1
X_15256_ _17329_/Q _09362_/C _15485_/B1 _16106_/Q vssd1 vssd1 vccd1 vccd1 _15256_/X
+ sky130_fd_sc_hd__a22o_1
X_12468_ _17327_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14207_ hold1533/X _14202_/B _14206_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14207_/X
+ sky130_fd_sc_hd__o211a_1
X_11419_ hold4941/X _12341_/B _11418_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11419_/X
+ sky130_fd_sc_hd__o211a_1
X_15187_ _15187_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15187_/X sky130_fd_sc_hd__or2_1
X_12399_ hold443/X hold589/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12400_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ hold735/X _14138_/B vssd1 vssd1 vccd1 vccd1 _14138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ hold2493/X _14105_/A2 _14068_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08630_ _13002_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _15937_/D sky130_fd_sc_hd__and2_1
X_17828_ _17862_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08561_ _09021_/A _08561_/B vssd1 vssd1 vccd1 vccd1 _15904_/D sky130_fd_sc_hd__and2_1
X_17759_ _17887_/CLK _17759_/D vssd1 vssd1 vccd1 vccd1 hold894/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_183_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18222_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08492_ _14330_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ hold2511/X _09119_/A2 _09112_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09044_ hold140/X hold659/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold420 hold420/A vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/A vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 input36/X vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold453 hold453/A vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold464 hold464/A vssd1 vssd1 vccd1 vccd1 input43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 hold486/A vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout900 _15187_/A vssd1 vssd1 vccd1 vccd1 _14740_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold497 data_in[13] vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 hold799/X vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__buf_4
XFILLER_0_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout922 hold729/X vssd1 vssd1 vccd1 vccd1 hold730/A sky130_fd_sc_hd__buf_4
XFILLER_0_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09946_ hold4198/X _10571_/B _09945_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09946_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout933 hold1452/X vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__buf_8
Xfanout944 hold746/X vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__buf_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ hold3463/X _10067_/B _09876_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09877_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _07795_/X vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _09149_/X vssd1 vssd1 vccd1 vccd1 _16187_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _15591_/Q vssd1 vssd1 vccd1 vccd1 hold1142/X sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ hold81/X _16033_/Q _08860_/S vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__mux2_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 _14829_/X vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _07998_/X vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _17925_/Q vssd1 vssd1 vccd1 vccd1 hold1175/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _09157_/X vssd1 vssd1 vccd1 vccd1 _16191_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ hold71/X hold632/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__mux2_1
Xhold1197 _17944_/Q vssd1 vssd1 vccd1 vccd1 hold1197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _12343_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__nor2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ hold932/X _16731_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ _13737_/A _13440_/B vssd1 vssd1 vccd1 vccd1 _13440_/X sky130_fd_sc_hd__or2_1
X_10652_ hold1956/X _16708_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ _13779_/A _13371_/B vssd1 vssd1 vccd1 vccd1 _13371_/X sky130_fd_sc_hd__or2_1
X_10583_ _16685_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__and3_1
XFILLER_0_146_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12322_ _13864_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _12322_/Y sky130_fd_sc_hd__nor2_1
X_15110_ hold863/X _15109_/B _15109_/Y _15032_/A vssd1 vssd1 vccd1 vccd1 hold864/A
+ sky130_fd_sc_hd__o211a_1
X_16090_ _17287_/CLK _16090_/D vssd1 vssd1 vccd1 vccd1 hold535/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ _14988_/A hold2262/X hold302/X vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ hold4997/X _12347_/B _12252_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ _11204_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__and3_1
X_12184_ hold4761/X _13844_/B _12183_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12184_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ hold2969/X _16869_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _11136_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16992_ _17893_/CLK _16992_/D vssd1 vssd1 vccd1 vccd1 _16992_/Q sky130_fd_sc_hd__dfxtp_1
X_15943_ _18406_/CLK _15943_/D vssd1 vssd1 vccd1 vccd1 hold592/A sky130_fd_sc_hd__dfxtp_1
X_11066_ hold1563/X hold5572/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__mux2_1
X_10017_ _13158_/A _09987_/A _10016_/X vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15874_ _17217_/CLK hold811/X vssd1 vssd1 vccd1 vccd1 hold810/A sky130_fd_sc_hd__dfxtp_1
X_17613_ _17741_/CLK _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14825_ hold1233/X _14828_/B _14824_/Y _14384_/A vssd1 vssd1 vccd1 vccd1 _14825_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _18360_/CLK _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _14988_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ hold4895/X _12347_/B _11967_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _13710_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__or2_1
X_17475_ _17475_/CLK _17475_/D vssd1 vssd1 vccd1 vccd1 _17475_/Q sky130_fd_sc_hd__dfxtp_1
X_10919_ hold1546/X _16797_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__mux2_1
X_11899_ hold4763/X _12377_/B _11898_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14687_ hold2803/X _14720_/B _14686_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14687_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ _18371_/CLK _16426_/D vssd1 vssd1 vccd1 vccd1 _16426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _13800_/A _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16357_ _18304_/CLK _16357_/D vssd1 vssd1 vccd1 vccd1 _16357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13569_ _13764_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13569_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ hold712/X _09386_/A _09392_/D hold560/X vssd1 vssd1 vccd1 vccd1 _15308_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5408 _10831_/X vssd1 vssd1 vccd1 vccd1 _16767_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16288_ _17511_/CLK _16288_/D vssd1 vssd1 vccd1 vccd1 _16288_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5419 _16463_/Q vssd1 vssd1 vccd1 vccd1 hold5419/X sky130_fd_sc_hd__dlygate4sd3_1
X_18027_ _18061_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15239_ hold426/X _15485_/A2 _15447_/B1 hold376/X _15238_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4707 _10210_/X vssd1 vssd1 vccd1 vccd1 _16560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4718 _17246_/Q vssd1 vssd1 vccd1 vccd1 hold4718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4729 _17220_/Q vssd1 vssd1 vccd1 vccd1 hold4729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout207 _11222_/B vssd1 vssd1 vccd1 vccd1 _11765_/B sky130_fd_sc_hd__buf_4
X_09800_ hold1091/X hold4319/X _11066_/S vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__mux2_1
Xfanout218 _10028_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__buf_4
X_07992_ hold606/A hold298/X hold624/A hold279/X vssd1 vssd1 vccd1 vccd1 _14681_/A
+ sky130_fd_sc_hd__nand4b_4
Xfanout229 _10610_/B vssd1 vssd1 vccd1 vccd1 _10897_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ hold485/X _16401_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09662_ hold1725/X _16378_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08613_ hold47/X hold268/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08614_/B sky130_fd_sc_hd__mux2_1
X_09593_ hold1373/X _13310_/A _10481_/S vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08544_ hold26/X hold519/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__mux2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08475_ hold5950/X _08486_/B _08474_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _08475_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17528_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09027_ _12422_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _16130_/D sky130_fd_sc_hd__and2_1
Xhold5920 _17550_/Q vssd1 vssd1 vccd1 vccd1 hold5920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5931 _17536_/Q vssd1 vssd1 vccd1 vccd1 hold5931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5942 hold6000/X vssd1 vssd1 vccd1 vccd1 hold5942/X sky130_fd_sc_hd__buf_1
Xhold5953 _15839_/Q vssd1 vssd1 vccd1 vccd1 hold5953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5964 _17948_/Q vssd1 vssd1 vccd1 vccd1 hold5964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 input21/X vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5975 _18335_/Q vssd1 vssd1 vccd1 vccd1 hold5975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5986 data_in[25] vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__clkbuf_4
Xhold5997 _18409_/Q vssd1 vssd1 vccd1 vccd1 hold5997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout730 _09011_/A vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__buf_2
Xfanout741 fanout763/X vssd1 vssd1 vccd1 vccd1 _13771_/C1 sky130_fd_sc_hd__buf_4
X_09929_ _18380_/Q hold4059/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__mux2_1
Xfanout752 _13909_/A vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__buf_4
Xfanout763 fanout842/X vssd1 vssd1 vccd1 vccd1 fanout763/X sky130_fd_sc_hd__buf_4
Xfanout774 _12274_/C1 vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__buf_4
Xfanout785 _14203_/C1 vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout796 fanout816/X vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ hold2451/X hold3587/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__mux2_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ hold2457/X hold3109/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12871_/X sky130_fd_sc_hd__mux2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _15105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_123 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _15219_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ hold2813/X _17098_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ _17274_/CLK _15590_/D vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _17075_/Q _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__and3_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14774_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__nand2_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11121_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__or2_1
X_17260_ _17260_/CLK _17260_/D vssd1 vssd1 vccd1 vccd1 _17260_/Q sky130_fd_sc_hd__dfxtp_1
X_11684_ _17900_/Q hold4601/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__mux2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ hold2717/X _14481_/B _14471_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _14472_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _17448_/CLK _16211_/D vssd1 vssd1 vccd1 vccd1 _16211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13423_ hold3504/X _13808_/B _13422_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13423_/X
+ sky130_fd_sc_hd__o211a_1
X_10635_ hold3630/X _10521_/A _10634_/X vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__a21oi_1
X_17191_ _18445_/CLK _17191_/D vssd1 vssd1 vccd1 vccd1 _17191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ _17329_/CLK _16142_/D vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13354_ hold4220/X _13832_/B _13353_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13354_/X
+ sky130_fd_sc_hd__o211a_1
X_10566_ hold3912/X _10563_/A _10565_/X vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12305_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12305_/X sky130_fd_sc_hd__and3_1
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16073_ _17345_/CLK _16073_/D vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__dfxtp_1
X_13285_ _13284_/X hold3728/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__mux2_1
X_10497_ _10521_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15024_ _15024_/A _15024_/B vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__and2_1
X_12236_ hold1216/X hold3444/X _12332_/C vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ hold2076/X hold4990/X _13388_/S vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _11121_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12098_ hold1457/X hold4024/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__mux2_1
X_16975_ _17887_/CLK _16975_/D vssd1 vssd1 vccd1 vccd1 _16975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15926_ _18405_/CLK _15926_/D vssd1 vssd1 vccd1 vccd1 hold419/A sky130_fd_sc_hd__dfxtp_1
X_11049_ _11637_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_0_127_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _17728_/CLK _15857_/D vssd1 vssd1 vccd1 vccd1 _15857_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14808_ hold883/X _14838_/B vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _17719_/CLK _15788_/D vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _17528_/CLK _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14739_ hold1557/X _14772_/B _14738_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14739_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08260_ _15539_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17458_ _18458_/CLK _17458_/D vssd1 vssd1 vccd1 vccd1 _17458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _18358_/CLK _16409_/D vssd1 vssd1 vccd1 vccd1 _16409_/Q sky130_fd_sc_hd__dfxtp_1
X_08191_ _15199_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _18441_/CLK _17389_/D vssd1 vssd1 vccd1 vccd1 _17389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5205 _17716_/Q vssd1 vssd1 vccd1 vccd1 hold5205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5216 _13765_/X vssd1 vssd1 vccd1 vccd1 _17708_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5227 _16916_/Q vssd1 vssd1 vccd1 vccd1 hold5227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5238 _11773_/Y vssd1 vssd1 vccd1 vccd1 _17081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4504 _17023_/Q vssd1 vssd1 vccd1 vccd1 hold4504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5249 _11217_/Y vssd1 vssd1 vccd1 vccd1 _11218_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4515 _11386_/X vssd1 vssd1 vccd1 vccd1 _16952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4526 _17701_/Q vssd1 vssd1 vccd1 vccd1 hold4526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4537 _12181_/X vssd1 vssd1 vccd1 vccd1 _17217_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3803 _10071_/Y vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4548 _10666_/X vssd1 vssd1 vccd1 vccd1 _16712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3814 _17582_/Q vssd1 vssd1 vccd1 vccd1 hold3814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4559 _17700_/Q vssd1 vssd1 vccd1 vccd1 hold4559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3825 _17103_/Q vssd1 vssd1 vccd1 vccd1 hold3825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3836 _12324_/Y vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3847 _13839_/Y vssd1 vssd1 vccd1 vccd1 _13840_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3858 _09907_/X vssd1 vssd1 vccd1 vccd1 _16459_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3869 _12348_/Y vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07975_ hold1816/X _07978_/B _07974_/Y _12831_/A vssd1 vssd1 vccd1 vccd1 _07975_/X
+ sky130_fd_sc_hd__o211a_1
X_09714_ _09948_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _09975_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__or2_1
X_09576_ _09954_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__or2_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _12422_/A hold510/X vssd1 vssd1 vccd1 vccd1 _15888_/D sky130_fd_sc_hd__and2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08458_ _15517_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08389_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ hold3338/X _10610_/B _10419_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10420_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ hold4317/X _10631_/B _10350_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13070_ _13070_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__or2_1
Xhold5750 _11113_/X vssd1 vssd1 vccd1 vccd1 _16861_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5761 hold5909/X vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__dlygate4sd3_1
X_10282_ hold5193/X _10628_/B _10281_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _10282_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5772 output87/X vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_12
Xhold5783 hold5918/X vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__dlygate4sd3_1
X_12021_ _13797_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5794 output91/X vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_286_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_215_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17829_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout560 _08173_/Y vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__clkbuf_8
Xfanout571 _07938_/Y vssd1 vssd1 vccd1 vccd1 _07991_/A2 sky130_fd_sc_hd__buf_6
Xfanout582 hold272/X vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__clkbuf_8
X_16760_ _18034_/CLK _16760_/D vssd1 vssd1 vccd1 vccd1 _16760_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout593 _12589_/S vssd1 vssd1 vccd1 vccd1 _12814_/S sky130_fd_sc_hd__clkbuf_8
X_13972_ _15207_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__or2_1
X_15711_ _17205_/CLK _15711_/D vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfxtp_1
X_12923_ hold3265/X _12922_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__mux2_1
X_16691_ _18217_/CLK _16691_/D vssd1 vssd1 vccd1 vccd1 _16691_/Q sky130_fd_sc_hd__dfxtp_1
X_18430_ _18450_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
X_15642_ _17282_/CLK _15642_/D vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ hold3199/X _12853_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__mux2_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _18395_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_11805_ _13797_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__or2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _17703_/CLK _15573_/D vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ hold3048/X _12784_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17331_/CLK _17312_/D vssd1 vssd1 vccd1 vccd1 hold387/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ hold2580/X _14541_/B _14523_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14524_/X
+ sky130_fd_sc_hd__o211a_1
X_18292_ _18324_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ hold3742/X _11640_/A _11735_/X vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17243_ _17275_/CLK _17243_/D vssd1 vssd1 vccd1 vccd1 _17243_/Q sky130_fd_sc_hd__dfxtp_1
X_14455_ _15189_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _11667_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ hold1146/X hold3185/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13407_/B sky130_fd_sc_hd__mux2_1
X_17174_ _17906_/CLK _17174_/D vssd1 vssd1 vccd1 vccd1 _17174_/Q sky130_fd_sc_hd__dfxtp_1
X_10618_ _11194_/A _10618_/B vssd1 vssd1 vccd1 vccd1 _10618_/Y sky130_fd_sc_hd__nor2_1
X_11598_ _11694_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__or2_1
X_14386_ _14390_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _17992_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ _17525_/CLK _16125_/D vssd1 vssd1 vccd1 vccd1 hold700/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13337_ hold1208/X _17566_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__mux2_1
X_10549_ hold4085/X _10643_/B _10548_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16056_ _17287_/CLK _16056_/D vssd1 vssd1 vccd1 vccd1 hold593/A sky130_fd_sc_hd__dfxtp_1
X_13268_ hold3601/X _13267_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__mux2_1
X_15007_ hold835/X _15006_/B _15006_/Y _15007_/C1 vssd1 vssd1 vccd1 vccd1 hold836/A
+ sky130_fd_sc_hd__o211a_1
X_12219_ _12285_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__or2_1
X_13199_ _13311_/A1 _13197_/X _13198_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13199_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2409 _18156_/Q vssd1 vssd1 vccd1 vccd1 hold2409/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1708 _18120_/Q vssd1 vssd1 vccd1 vccd1 hold1708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 _15226_/X vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16958_ _17870_/CLK _16958_/D vssd1 vssd1 vccd1 vccd1 _16958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _17307_/CLK _15909_/D vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_16889_ _18033_/CLK _16889_/D vssd1 vssd1 vccd1 vccd1 _16889_/Q sky130_fd_sc_hd__dfxtp_1
X_09430_ hold616/X _16301_/Q vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09400_/A _09364_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__nor3_1
X_08312_ hold5978/X _08323_/B _08311_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08312_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ hold2644/X _09338_/A2 _09291_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_12 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_23 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ hold2842/X _08262_/B _08242_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08243_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_34 _15215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_5_31__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_31__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_56 _15535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 hold490/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _08504_/A _15182_/A vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__or2_4
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_78 hold883/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 hold5839/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5002 _12190_/X vssd1 vssd1 vccd1 vccd1 _17220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5013 _16583_/Q vssd1 vssd1 vccd1 vccd1 hold5013/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5024 _12067_/X vssd1 vssd1 vccd1 vccd1 _17179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5035 _12121_/X vssd1 vssd1 vccd1 vccd1 _17197_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5046 _17241_/Q vssd1 vssd1 vccd1 vccd1 hold5046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4301 _16834_/Q vssd1 vssd1 vccd1 vccd1 hold4301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4312 _11812_/X vssd1 vssd1 vccd1 vccd1 _17094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5057 _09562_/X vssd1 vssd1 vccd1 vccd1 _16344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4323 _16438_/Q vssd1 vssd1 vccd1 vccd1 hold4323/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput130 hold5869/X vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_12
Xhold5068 _17274_/Q vssd1 vssd1 vccd1 vccd1 hold5068/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput141 _13043_/C vssd1 vssd1 vccd1 vccd1 load_status[1] sky130_fd_sc_hd__buf_12
Xhold4334 _13615_/X vssd1 vssd1 vccd1 vccd1 _17658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5079 _12166_/X vssd1 vssd1 vccd1 vccd1 _17212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3600 _10003_/Y vssd1 vssd1 vccd1 vccd1 _16491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4345 _17699_/Q vssd1 vssd1 vccd1 vccd1 hold4345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4356 _11629_/X vssd1 vssd1 vccd1 vccd1 _17033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3611 _11142_/Y vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3622 _17565_/Q vssd1 vssd1 vccd1 vccd1 hold3622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4367 _17001_/Q vssd1 vssd1 vccd1 vccd1 hold4367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3633 _16524_/Q vssd1 vssd1 vccd1 vccd1 hold3633/X sky130_fd_sc_hd__buf_2
Xhold4378 _13384_/X vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4389 _17154_/Q vssd1 vssd1 vccd1 vccd1 hold4389/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3644 _10645_/Y vssd1 vssd1 vccd1 vccd1 _16705_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2910 _14175_/X vssd1 vssd1 vccd1 vccd1 _17890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3655 _10035_/Y vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3666 _11160_/Y vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2921 _18020_/Q vssd1 vssd1 vccd1 vccd1 hold2921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2932 _18325_/Q vssd1 vssd1 vccd1 vccd1 hold2932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3677 _10060_/Y vssd1 vssd1 vccd1 vccd1 _16510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3688 _13821_/Y vssd1 vssd1 vccd1 vccd1 _13822_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 _18377_/Q vssd1 vssd1 vccd1 vccd1 hold2943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2954 _09131_/X vssd1 vssd1 vccd1 vccd1 _16178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3699 _16546_/Q vssd1 vssd1 vccd1 vccd1 hold3699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2965 _18351_/Q vssd1 vssd1 vccd1 vccd1 hold2965/X sky130_fd_sc_hd__dlygate4sd3_1
X_07958_ _15527_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07958_/X sky130_fd_sc_hd__or2_1
Xhold2976 _14061_/X vssd1 vssd1 vccd1 vccd1 _17835_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2987 _15726_/Q vssd1 vssd1 vccd1 vccd1 hold2987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 _08290_/X vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07889_ hold1126/X _07918_/B _07888_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _07889_/X
+ sky130_fd_sc_hd__o211a_1
X_09628_ hold3861/X _10028_/B _09627_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ hold3562/X _10049_/B _09558_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09559_/X
+ sky130_fd_sc_hd__o211a_1
X_12570_ _12996_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _17366_/D sky130_fd_sc_hd__and2_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11521_ hold4686/X _12305_/B _11520_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11521_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11452_ hold4419/X _11735_/B _11451_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11452_/X
+ sky130_fd_sc_hd__o211a_1
X_14240_ _15189_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ hold2799/X _16625_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10404_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14171_ hold1661/X _14198_/B _14170_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _14171_/X
+ sky130_fd_sc_hd__o211a_1
X_11383_ hold5715/X _11765_/B _11382_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10334_ hold1557/X hold4242/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _17566_/Q _17100_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13053_ _13053_/A _13056_/C _13055_/C _13046_/A vssd1 vssd1 vccd1 vccd1 _13230_/B
+ sky130_fd_sc_hd__or4b_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5580 _16979_/Q vssd1 vssd1 vccd1 vccd1 hold5580/X sky130_fd_sc_hd__dlygate4sd3_1
X_17930_ _18158_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
X_10265_ hold1436/X hold3206/X _10649_/C vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5591 _11137_/X vssd1 vssd1 vccd1 vccd1 _16869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12004_ hold4024/X _13811_/B _12003_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12004_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4890 _13516_/X vssd1 vssd1 vccd1 vccd1 _17625_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17861_ _17873_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
X_10196_ hold1473/X _16556_/Q _10643_/C vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _18461_/CLK _16812_/D vssd1 vssd1 vccd1 vccd1 _16812_/Q sky130_fd_sc_hd__dfxtp_1
X_17792_ _17855_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout390 _14718_/B vssd1 vssd1 vccd1 vccd1 _14720_/B sky130_fd_sc_hd__buf_6
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16743_ _18043_/CLK _16743_/D vssd1 vssd1 vccd1 vccd1 _16743_/Q sky130_fd_sc_hd__dfxtp_1
X_13955_ hold1679/X _13980_/B _13954_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _13955_/X
+ sky130_fd_sc_hd__o211a_1
X_12906_ _12909_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _17478_/D sky130_fd_sc_hd__and2_1
X_16674_ _18224_/CLK _16674_/D vssd1 vssd1 vccd1 vccd1 _16674_/Q sky130_fd_sc_hd__dfxtp_1
X_13886_ _17749_/Q _13886_/B _13886_/C vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__and3_1
X_18413_ _18413_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15625_ _17221_/CLK _15625_/D vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12843_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _17455_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18381_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15556_ hold2734/X _15560_/A2 _15555_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _15556_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12768_ _12804_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _17432_/D sky130_fd_sc_hd__and2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ _14972_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11719_ _12301_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11719_/Y sky130_fd_sc_hd__nor2_1
X_18275_ _18371_/CLK hold953/X vssd1 vssd1 vccd1 vccd1 hold952/A sky130_fd_sc_hd__dfxtp_1
X_15487_ _17324_/Q _09357_/A _15487_/B1 hold620/X _15486_/X vssd1 vssd1 vccd1 vccd1
+ _15489_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ _12789_/A _12699_/B vssd1 vssd1 vccd1 vccd1 _17409_/D sky130_fd_sc_hd__and2_1
X_17226_ _18445_/CLK _17226_/D vssd1 vssd1 vccd1 vccd1 _17226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 input10/A vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14438_ hold1154/X hold209/X _14437_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _14438_/X
+ sky130_fd_sc_hd__o211a_1
Xinput21 input21/A vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput32 input32/A vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput43 input43/A vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
Xinput54 input54/A vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
X_17157_ _17221_/CLK _17157_/D vssd1 vssd1 vccd1 vccd1 _17157_/Q sky130_fd_sc_hd__dfxtp_1
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
Xhold805 hold805/A vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _15103_/A hold2167/X hold275/X vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_137_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18360_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16108_ _17331_/CLK _16108_/D vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__dfxtp_1
Xhold827 hold827/A vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 hold838/A vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 la_data_in[25] vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _17893_/CLK _17088_/D vssd1 vssd1 vccd1 vccd1 _17088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16039_ _18415_/CLK _16039_/D vssd1 vssd1 vccd1 vccd1 hold595/A sky130_fd_sc_hd__dfxtp_1
X_08930_ hold14/X hold532/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08931_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2206 _09231_/X vssd1 vssd1 vccd1 vccd1 _16227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 _08214_/X vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08861_ _15454_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _16049_/D sky130_fd_sc_hd__and2_1
Xhold2228 _16192_/Q vssd1 vssd1 vccd1 vccd1 hold2228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2239 _15658_/Q vssd1 vssd1 vccd1 vccd1 hold2239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 _18102_/Q vssd1 vssd1 vccd1 vccd1 hold1505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 _14685_/X vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ _16286_/Q _07810_/Y hold1772/X _09339_/B vssd1 vssd1 vccd1 vccd1 _07812_/Y
+ sky130_fd_sc_hd__a31oi_1
X_08792_ _15473_/A _08792_/B vssd1 vssd1 vccd1 vccd1 _16016_/D sky130_fd_sc_hd__and2_1
Xhold1527 _18259_/Q vssd1 vssd1 vccd1 vccd1 hold1527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _18154_/Q vssd1 vssd1 vccd1 vccd1 hold1538/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 _07983_/X vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _07804_/A _09456_/C _15334_/A _09412_/X vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ _15543_/A hold265/A _15182_/A _09352_/D vssd1 vssd1 vccd1 vccd1 _09363_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09275_ _15551_/A hold1407/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08226_ hold1990/X _08209_/B _08225_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08157_ _08504_/A _15492_/A vssd1 vssd1 vccd1 vccd1 _08170_/S sky130_fd_sc_hd__nand2b_4
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08088_ _14774_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4120 _10819_/X vssd1 vssd1 vccd1 vccd1 _16763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4131 _16751_/Q vssd1 vssd1 vccd1 vccd1 hold4131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4142 _10297_/X vssd1 vssd1 vccd1 vccd1 _16589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4153 _16994_/Q vssd1 vssd1 vccd1 vccd1 hold4153/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4164 _13438_/X vssd1 vssd1 vccd1 vccd1 _17599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4175 _10546_/X vssd1 vssd1 vccd1 vccd1 _16672_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3430 _12938_/X vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10050_ _13246_/A _09954_/A _10049_/X vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__a21oi_1
Xhold3441 _11494_/X vssd1 vssd1 vccd1 vccd1 _16988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4186 _16827_/Q vssd1 vssd1 vccd1 vccd1 hold4186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4197 _10393_/X vssd1 vssd1 vccd1 vccd1 _16621_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3452 _12995_/X vssd1 vssd1 vccd1 vccd1 _12996_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3463 _16481_/Q vssd1 vssd1 vccd1 vccd1 hold3463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3474 _17165_/Q vssd1 vssd1 vccd1 vccd1 hold3474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3485 _09589_/X vssd1 vssd1 vccd1 vccd1 _16353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2740 _17958_/Q vssd1 vssd1 vccd1 vccd1 hold2740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2751 _09229_/X vssd1 vssd1 vccd1 vccd1 _16226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3496 _11944_/X vssd1 vssd1 vccd1 vccd1 _17138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2762 _17887_/Q vssd1 vssd1 vccd1 vccd1 hold2762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2773 _08241_/X vssd1 vssd1 vccd1 vccd1 _15755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2784 _14177_/X vssd1 vssd1 vccd1 vccd1 _17891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2795 _15860_/Q vssd1 vssd1 vccd1 vccd1 hold2795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _13776_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13740_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ hold1306/X _16808_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13671_ _13767_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__or2_1
X_10883_ hold483/X hold3275/X _11747_/C vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__mux2_1
X_15410_ hold419/X _15486_/A2 _15446_/B1 hold461/X vssd1 vssd1 vccd1 vccd1 _15410_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12622_ hold1529/X _17385_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__mux2_1
X_16390_ _18337_/CLK _16390_/D vssd1 vssd1 vccd1 vccd1 _16390_/Q sky130_fd_sc_hd__dfxtp_1
X_15341_ _16298_/Q _15477_/A2 _15487_/B1 hold396/X _15340_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ hold2566/X hold3244/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11504_ hold1082/X _16992_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__mux2_1
X_18060_ _18060_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15272_ _15489_/A _15272_/B _15272_/C _15272_/D vssd1 vssd1 vccd1 vccd1 _15272_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _17335_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__or2_1
X_17011_ _17891_/CLK _17011_/D vssd1 vssd1 vccd1 vccd1 _17011_/Q sky130_fd_sc_hd__dfxtp_1
X_14223_ hold1979/X _14216_/Y _14222_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11435_ hold2004/X _16969_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_230_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14154_ _15553_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14154_/X sky130_fd_sc_hd__or2_1
X_11366_ hold1744/X _16946_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ _13105_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__and2_1
X_10317_ _10527_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _17771_/Q hold3781/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__mux2_1
X_14085_ hold2330/X _14094_/B _14084_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14085_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13053_/A _13035_/X hold901/X vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__mux2_1
X_10248_ _10542_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__or2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _18072_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17844_ _17844_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10179_ _10563_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10179_/X sky130_fd_sc_hd__or2_1
X_17775_ _18032_/CLK hold732/X vssd1 vssd1 vccd1 vccd1 _17775_/Q sky130_fd_sc_hd__dfxtp_1
X_14987_ hold2487/X _15004_/B _14986_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _14987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16726_ _18059_/CLK _16726_/D vssd1 vssd1 vccd1 vccd1 _16726_/Q sky130_fd_sc_hd__dfxtp_1
X_13938_ _14726_/A hold1919/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _18215_/CLK _16657_/D vssd1 vssd1 vccd1 vccd1 _16657_/Q sky130_fd_sc_hd__dfxtp_1
X_13869_ hold3822/X _13776_/A _13868_/X vssd1 vssd1 vccd1 vccd1 _13869_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15608_ _17453_/CLK _15608_/D vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _18210_/CLK _16588_/D vssd1 vssd1 vccd1 vccd1 _16588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18327_ _18353_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15539_ _15539_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09060_ hold14/X hold445/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__mux2_1
X_18258_ _18358_/CLK hold832/X vssd1 vssd1 vccd1 vccd1 hold831/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_318_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17691_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ _15525_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__or2_1
X_17209_ _17703_/CLK _17209_/D vssd1 vssd1 vccd1 vccd1 _17209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _18221_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold602 hold602/A vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 hold613/A vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 hold624/A vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold635 hold635/A vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 hold646/A vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 hold657/A vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold668 hold668/A vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 hold679/A vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ hold2002/X hold5588/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ _15284_/A _08913_/B vssd1 vssd1 vccd1 vccd1 _16074_/D sky130_fd_sc_hd__and2_1
Xhold2003 _15218_/X vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09893_ hold2078/X _16455_/Q _09893_/S vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__mux2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2014 _15649_/Q vssd1 vssd1 vccd1 vccd1 hold2014/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _08281_/X vssd1 vssd1 vccd1 vccd1 _15775_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2036 _18021_/Q vssd1 vssd1 vccd1 vccd1 hold2036/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _15884_/Q vssd1 vssd1 vccd1 vccd1 hold1302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2047 _14269_/X vssd1 vssd1 vccd1 vccd1 _17935_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ hold5/X hold470/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__mux2_1
Xhold1313 _18437_/Q vssd1 vssd1 vccd1 vccd1 hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2058 _18342_/Q vssd1 vssd1 vccd1 vccd1 hold2058/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 _18213_/Q vssd1 vssd1 vccd1 vccd1 hold1324/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _14482_/X vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 _15754_/Q vssd1 vssd1 vccd1 vccd1 hold1335/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1346 _18444_/Q vssd1 vssd1 vccd1 vccd1 hold1346/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1357 _17807_/Q vssd1 vssd1 vccd1 vccd1 hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _18294_/Q vssd1 vssd1 vccd1 vccd1 hold1368/X sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ hold140/X _16008_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__mux2_1
Xhold1379 _18245_/Q vssd1 vssd1 vccd1 vccd1 hold1379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18009_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _15169_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _12756_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _16240_/D sky130_fd_sc_hd__and2_1
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08209_ _15217_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09189_ hold1179/X _09216_/B _09188_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _09189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11220_ hold3705/X _11031_/A _11219_/X vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11151_ hold3616/X _11061_/A _11150_/X vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ hold4190/X _10580_/B _10101_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10102_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11082_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3260 _17472_/Q vssd1 vssd1 vccd1 vccd1 hold3260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3271 _16671_/Q vssd1 vssd1 vccd1 vccd1 hold3271/X sky130_fd_sc_hd__dlygate4sd3_1
X_10033_ _10588_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10033_/Y sky130_fd_sc_hd__nor2_1
X_14910_ _14980_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3282 _17475_/Q vssd1 vssd1 vccd1 vccd1 hold3282/X sky130_fd_sc_hd__dlygate4sd3_1
X_15890_ _18409_/CLK _15890_/D vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__dfxtp_1
Xhold3293 _17598_/Q vssd1 vssd1 vccd1 vccd1 hold3293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2570 _18234_/Q vssd1 vssd1 vccd1 vccd1 hold2570/X sky130_fd_sc_hd__dlygate4sd3_1
X_14841_ hold2266/X _14828_/B _14840_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14841_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2581 _14524_/X vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2592 _18104_/Q vssd1 vssd1 vccd1 vccd1 hold2592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ _17725_/CLK _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1880 _09219_/X vssd1 vssd1 vccd1 vccd1 _16221_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14772_ _15219_/A _14772_/B vssd1 vssd1 vccd1 vccd1 _14772_/Y sky130_fd_sc_hd__nand2_1
Xhold1891 _15734_/Q vssd1 vssd1 vccd1 vccd1 hold1891/X sky130_fd_sc_hd__dlygate4sd3_1
X_11984_ hold1163/X hold3315/X _12368_/C vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__mux2_1
X_16511_ _18185_/CLK _16511_/D vssd1 vssd1 vccd1 vccd1 _16511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13723_ hold4411/X _13862_/B _13722_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__o211a_1
X_10935_ _11694_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17491_ _17494_/CLK _17491_/D vssd1 vssd1 vccd1 vccd1 _17491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16442_ _18355_/CLK _16442_/D vssd1 vssd1 vccd1 vccd1 _16442_/Q sky130_fd_sc_hd__dfxtp_1
X_13654_ hold3566/X _13886_/B _13653_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _11067_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ hold3257/X _12604_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__mux2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _18382_/CLK _16373_/D vssd1 vssd1 vccd1 vccd1 _16373_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ hold4673/X _13868_/B _13584_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10797_ _11097_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__or2_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18112_ _18176_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15324_ _15414_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__and2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ hold3597/X _12535_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _18043_/CLK hold575/X vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ hold452/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12467_ hold53/X _12445_/A _12505_/A3 _12466_/X _15491_/A vssd1 vssd1 vccd1 vccd1
+ hold54/A sky130_fd_sc_hd__o311a_1
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _14330_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14206_/X sky130_fd_sc_hd__or2_1
X_11418_ _12246_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__or2_1
X_15186_ hold1363/X _15219_/B _15185_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _15186_/X
+ sky130_fd_sc_hd__o211a_1
X_12398_ _12438_/A _12398_/B vssd1 vssd1 vccd1 vccd1 _17292_/D sky130_fd_sc_hd__and2_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ hold1734/X hold587/X _14136_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14137_/X
+ sky130_fd_sc_hd__o211a_1
X_11349_ _12018_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__or2_1
X_14068_ _14246_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14068_/X sky130_fd_sc_hd__or2_1
X_13019_ hold925/X input1/X hold898/X hold792/X vssd1 vssd1 vccd1 vccd1 hold926/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17827_ _17827_/CLK hold842/X vssd1 vssd1 vccd1 vccd1 hold841/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ hold71/X hold349/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08561_/B sky130_fd_sc_hd__mux2_1
X_17758_ _17923_/CLK _17758_/D vssd1 vssd1 vccd1 vccd1 _17758_/Q sky130_fd_sc_hd__dfxtp_1
X_08491_ hold810/X _08486_/B _08490_/X _08149_/A vssd1 vssd1 vccd1 vccd1 hold811/A
+ sky130_fd_sc_hd__o211a_1
X_16709_ _18042_/CLK _16709_/D vssd1 vssd1 vccd1 vccd1 _16709_/Q sky130_fd_sc_hd__dfxtp_1
X_17689_ _17721_/CLK _17689_/D vssd1 vssd1 vccd1 vccd1 _17689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09112_ _15553_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_152_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18197_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09043_ _15304_/A _09043_/B vssd1 vssd1 vccd1 vccd1 _16138_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold410 data_in[17] vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/A vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold443/A vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__buf_4
Xhold454 hold454/A vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 input43/X vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__buf_1
Xhold476 hold476/A vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 hold58/X vssd1 vssd1 vccd1 vccd1 input9/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 hold1057/X vssd1 vssd1 vccd1 vccd1 hold1058/A sky130_fd_sc_hd__buf_6
Xfanout912 hold798/X vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__buf_6
X_09945_ _10380_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__or2_1
Xfanout923 hold891/X vssd1 vssd1 vccd1 vccd1 hold892/A sky130_fd_sc_hd__buf_6
Xfanout934 hold1452/X vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__buf_8
Xfanout945 hold944/X vssd1 vssd1 vccd1 vccd1 _14218_/A sky130_fd_sc_hd__buf_6
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09951_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__or2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _18200_/Q vssd1 vssd1 vccd1 vccd1 hold1110/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _07796_/Y vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _17828_/Q vssd1 vssd1 vccd1 vccd1 hold1132/X sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _12438_/A hold166/X vssd1 vssd1 vccd1 vccd1 _16032_/D sky130_fd_sc_hd__and2_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _07895_/X vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1154 _18017_/Q vssd1 vssd1 vccd1 vccd1 hold1154/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _17792_/Q vssd1 vssd1 vccd1 vccd1 hold1165/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 _14249_/X vssd1 vssd1 vccd1 vccd1 _17925_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _15835_/Q vssd1 vssd1 vccd1 vccd1 hold1187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _15304_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _15999_/D sky130_fd_sc_hd__and2_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _14289_/X vssd1 vssd1 vccd1 vccd1 _17944_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ hold81/X hold549/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__mux2_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ hold5574/X _11213_/B _10719_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10720_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ _11194_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10582_/Y sky130_fd_sc_hd__nor2_1
X_13370_ _15866_/Q hold3919/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13371_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ hold3805/X _12093_/A _12320_/X vssd1 vssd1 vccd1 vccd1 _12321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15040_ _15044_/A _15040_/B vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__and2_1
X_12252_ _12255_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__or2_1
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_181_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12183_ _13749_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
X_11134_ hold4149/X _11735_/B _11133_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11134_/X
+ sky130_fd_sc_hd__o211a_1
X_16991_ _17903_/CLK _16991_/D vssd1 vssd1 vccd1 vccd1 _16991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15942_ _17289_/CLK _15942_/D vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__dfxtp_1
X_11065_ hold5649/X _09992_/B _11064_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _11065_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3090 _12683_/X vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10016_ _16496_/Q _10016_/B _10022_/C vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__and3_1
X_15873_ _17742_/CLK _15873_/D vssd1 vssd1 vccd1 vccd1 _15873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17612_ _17740_/CLK _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_1
X_14824_ _15109_/A _14828_/B vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _18360_/CLK _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ hold2612/X _14772_/B _14754_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14755_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _12255_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__or2_1
XFILLER_0_169_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ hold1987/X hold4775/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__mux2_1
X_17474_ _17475_/CLK _17474_/D vssd1 vssd1 vccd1 vccd1 _17474_/Q sky130_fd_sc_hd__dfxtp_1
X_10918_ hold3886/X _11210_/B _10917_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14686_ _14740_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11898_ _12282_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__or2_1
X_16425_ _18415_/CLK _16425_/D vssd1 vssd1 vccd1 vccd1 _16425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13637_ hold2464/X hold4463/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ hold5468/X _11156_/B _10848_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ _18397_/CLK _16356_/D vssd1 vssd1 vccd1 vccd1 _16356_/Q sky130_fd_sc_hd__dfxtp_1
X_13568_ hold1242/X hold4595/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ hold659/X _15479_/A2 _09386_/D hold536/X _15306_/X vssd1 vssd1 vccd1 vccd1
+ _15312_/B sky130_fd_sc_hd__a221o_1
X_12519_ _13002_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _17349_/D sky130_fd_sc_hd__and2_1
XFILLER_0_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16287_ _18462_/CLK _16287_/D vssd1 vssd1 vccd1 vccd1 _16287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13499_ hold1669/X _17620_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13500_/B sky130_fd_sc_hd__mux2_1
Xhold5409 _16980_/Q vssd1 vssd1 vccd1 vccd1 hold5409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18026_ _18067_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15238_ hold418/X _15484_/A2 _15451_/A2 hold475/X vssd1 vssd1 vccd1 vccd1 _15238_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4708 _17735_/Q vssd1 vssd1 vccd1 vccd1 hold4708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4719 _12172_/X vssd1 vssd1 vccd1 vccd1 _17214_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15169_ _15169_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15169_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout208 fanout209/X vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__buf_4
Xfanout219 _09517_/A2 vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07991_ hold2133/X _07991_/A2 _07990_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _07991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ hold5643/X _11201_/B _09729_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _09730_/X
+ sky130_fd_sc_hd__o211a_1
X_09661_ hold4279/X _10049_/B _09660_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09661_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08612_ _09021_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _15928_/D sky130_fd_sc_hd__and2_1
X_09592_ hold4692/X _10070_/B _09591_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09592_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _09003_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _15895_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ _15207_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5910 _17543_/Q vssd1 vssd1 vccd1 vccd1 hold5910/X sky130_fd_sc_hd__dlygate4sd3_1
X_09026_ hold59/X hold591/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5921 _17538_/Q vssd1 vssd1 vccd1 vccd1 hold5921/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5932 _17557_/Q vssd1 vssd1 vccd1 vccd1 hold5932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5943 hold5999/X vssd1 vssd1 vccd1 vccd1 hold5943/X sky130_fd_sc_hd__buf_1
Xhold5954 _18240_/Q vssd1 vssd1 vccd1 vccd1 hold5954/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 hold652/X vssd1 vssd1 vccd1 vccd1 hold653/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5965 _17856_/Q vssd1 vssd1 vccd1 vccd1 hold5965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__clkbuf_4
Xhold5976 _18343_/Q vssd1 vssd1 vccd1 vccd1 hold5976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5987 data_in[26] vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 la_data_in[16] vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5998 data_in[31] vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold22/X vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 la_data_in[29] vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout720 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _15172_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout731 _08585_/A vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__buf_2
X_09928_ hold5631/X _10016_/B _09927_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09928_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout742 _08111_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__buf_4
Xfanout753 fanout763/X vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__buf_2
Xfanout764 _13753_/C1 vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__buf_4
Xfanout775 _12274_/C1 vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__buf_2
Xfanout786 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _14203_/C1 sky130_fd_sc_hd__clkbuf_4
X_09859_ hold4549/X _10049_/B _09858_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09859_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout797 _15072_/A vssd1 vssd1 vccd1 vccd1 _15007_/C1 sky130_fd_sc_hd__buf_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12924_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _17466_/D sky130_fd_sc_hd__and2_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _15103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ hold4769/X _12299_/B _11820_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11821_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ hold2641/X _14541_/B _14539_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14540_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _12331_/A _11752_/B vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__nor2_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ hold2485/X hold5251/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__mux2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _15205_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14471_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11683_ hold4621/X _12323_/B _11682_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11683_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16210_ _17448_/CLK _16210_/D vssd1 vssd1 vccd1 vccd1 _16210_/Q sky130_fd_sc_hd__dfxtp_1
X_13422_ _13713_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17190_ _17592_/CLK _17190_/D vssd1 vssd1 vccd1 vccd1 _17190_/Q sky130_fd_sc_hd__dfxtp_1
X_10634_ _16702_/Q _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10634_/X sky130_fd_sc_hd__and3_1
XFILLER_0_181_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _18409_/CLK _16141_/D vssd1 vssd1 vccd1 vccd1 hold375/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13353_ _13737_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ _16679_/Q _10568_/B _10565_/C vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__and3_1
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _13822_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12304_/Y sky130_fd_sc_hd__nor2_1
X_16072_ _17318_/CLK _16072_/D vssd1 vssd1 vccd1 vccd1 hold371/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13284_ hold5248/X _13283_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__mux2_1
X_10496_ hold1746/X hold4213/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__mux2_1
X_15023_ _15185_/A hold1614/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15024_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12235_ hold5522/X _12329_/B _12234_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _12235_/X
+ sky130_fd_sc_hd__o211a_1
X_12166_ hold5078/X _12356_/B _12165_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ hold2641/X _16863_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__mux2_1
X_12097_ hold4184/X _12308_/B _12096_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12097_/X
+ sky130_fd_sc_hd__o211a_1
X_16974_ _18051_/CLK _16974_/D vssd1 vssd1 vccd1 vccd1 _16974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15925_ _18413_/CLK _15925_/D vssd1 vssd1 vccd1 vccd1 hold548/A sky130_fd_sc_hd__dfxtp_1
X_11048_ _18043_/Q hold4451/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__mux2_1
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15856_ _17726_/CLK _15856_/D vssd1 vssd1 vccd1 vccd1 _15856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14807_ hold2774/X _14828_/B _14806_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14807_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15787_ _17686_/CLK _15787_/D vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _13002_/A _12999_/B vssd1 vssd1 vccd1 vccd1 _17509_/D sky130_fd_sc_hd__and2_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17526_ _18308_/CLK _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_1
X_14738_ _15185_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14738_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17457_ _18458_/CLK _17457_/D vssd1 vssd1 vccd1 vccd1 _17457_/Q sky130_fd_sc_hd__dfxtp_1
X_14669_ hold2115/X _14664_/B _14668_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _14669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_5_30__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_30__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_16408_ _18353_/CLK _16408_/D vssd1 vssd1 vccd1 vccd1 _16408_/Q sky130_fd_sc_hd__dfxtp_1
X_08190_ hold1426/X _08209_/B _08189_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ _18454_/CLK _17388_/D vssd1 vssd1 vccd1 vccd1 _17388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ _18386_/CLK _16339_/D vssd1 vssd1 vccd1 vccd1 _16339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5206 _13693_/X vssd1 vssd1 vccd1 vccd1 _17684_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5217 _16013_/Q vssd1 vssd1 vccd1 vccd1 _15435_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5228 _11757_/Y vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5239 _17107_/Q vssd1 vssd1 vccd1 vccd1 hold5239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4505 _11503_/X vssd1 vssd1 vccd1 vccd1 _16991_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4516 _16595_/Q vssd1 vssd1 vccd1 vccd1 hold4516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18009_ _18009_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4527 _13648_/X vssd1 vssd1 vccd1 vccd1 _17669_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4538 _17051_/Q vssd1 vssd1 vccd1 vccd1 hold4538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4549 _16475_/Q vssd1 vssd1 vccd1 vccd1 hold4549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3804 _10072_/Y vssd1 vssd1 vccd1 vccd1 _16514_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3815 _13866_/Y vssd1 vssd1 vccd1 vccd1 _13867_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3826 _12318_/Y vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3837 _12325_/Y vssd1 vssd1 vccd1 vccd1 _17265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3848 _13840_/Y vssd1 vssd1 vccd1 vccd1 _17733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3859 _16365_/Q vssd1 vssd1 vccd1 vccd1 hold3859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07974_ _15543_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07974_/Y sky130_fd_sc_hd__nand2_1
X_09713_ hold2643/X _16395_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ hold1385/X _16372_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09575_ hold1103/X _13262_/A _10055_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ hold68/X hold509/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold510/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ hold1644/X _08488_/B _08456_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _08457_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08388_ _15123_/A _15826_/Q _08390_/S vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _10524_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _12438_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _16121_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5740 _11290_/X vssd1 vssd1 vccd1 vccd1 _16920_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5751 hold5904/X vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__buf_1
X_10281_ _10491_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5762 output81/X vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_12
XFILLER_0_143_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5773 hold5915/X vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5784 hold5784/A vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_12
X_12020_ hold1606/X hold3242/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__mux2_1
Xhold5795 hold5926/X vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout550 hold121/X vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__buf_6
Xfanout561 hold195/X vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__buf_6
Xfanout572 _07916_/B vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__buf_6
Xfanout583 _13057_/X vssd1 vssd1 vccd1 vccd1 _13250_/S sky130_fd_sc_hd__buf_8
X_13971_ hold1165/X _13980_/B _13970_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _13971_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout594 _12679_/S vssd1 vssd1 vccd1 vccd1 _12844_/S sky130_fd_sc_hd__clkbuf_8
X_15710_ _17584_/CLK hold198/X vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_255_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12922_ hold2121/X _17485_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux2_1
X_16690_ _18216_/CLK _16690_/D vssd1 vssd1 vccd1 vccd1 _16690_/Q sky130_fd_sc_hd__dfxtp_1
X_15641_ _17279_/CLK _15641_/D vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfxtp_1
X_12853_ hold2953/X _17462_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__mux2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18360_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
X_11804_ hold2396/X hold4925/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__mux2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15572_ _17906_/CLK _15572_/D vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ hold2376/X _17439_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__mux2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _18421_/CLK _17311_/D vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__dfxtp_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14988_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__or2_1
X_18291_ _18324_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11735_ _17069_/Q _11735_/B _11735_/C vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__and3_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17274_/CLK _17242_/D vssd1 vssd1 vccd1 vccd1 _17242_/Q sky130_fd_sc_hd__dfxtp_1
X_14454_ hold2878/X _14481_/B _14453_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _14454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ hold1084/X _17046_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ hold5213/X _13883_/B _13404_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17173_ _17779_/CLK _17173_/D vssd1 vssd1 vccd1 vccd1 _17173_/Q sky130_fd_sc_hd__dfxtp_1
X_10617_ hold3619/X _10521_/A _10616_/X vssd1 vssd1 vccd1 vccd1 _10617_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14385_ _14726_/A hold1849/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ hold1491/X hold4504/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16124_ _17531_/CLK _16124_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
X_13336_ hold4496/X _13814_/B _13335_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13336_/X
+ sky130_fd_sc_hd__o211a_1
X_10548_ _10548_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16055_ _18409_/CLK _16055_/D vssd1 vssd1 vccd1 vccd1 hold454/A sky130_fd_sc_hd__dfxtp_1
X_13267_ _13266_/X _16926_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__mux2_1
X_10479_ _11082_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15006_ _15221_/A _15006_/B vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nand2_1
X_12218_ hold1094/X _17230_/Q _12353_/C vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__mux2_1
X_13198_ _13198_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ hold1142/X hold4593/X _12377_/C vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1709 _14655_/X vssd1 vssd1 vccd1 vccd1 _18120_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16957_ _17892_/CLK _16957_/D vssd1 vssd1 vccd1 vccd1 _16957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15908_ _18425_/CLK _15908_/D vssd1 vssd1 vccd1 vccd1 hold715/A sky130_fd_sc_hd__dfxtp_1
X_16888_ _18228_/CLK _16888_/D vssd1 vssd1 vccd1 vccd1 _16888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15839_ _17634_/CLK _15839_/D vssd1 vssd1 vccd1 vccd1 _15839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _09400_/A _09360_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09360_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08311_ _08311_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__or2_1
X_17509_ _17517_/CLK _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09291_ _14972_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _13164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ _14246_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08242_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_24 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _15215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_46 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _14866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17511_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_68 hold667/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08173_ _08504_/A _15182_/A vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_79 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5003 _16962_/Q vssd1 vssd1 vccd1 vccd1 hold5003/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5014 _10183_/X vssd1 vssd1 vccd1 vccd1 _16551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5025 _17590_/Q vssd1 vssd1 vccd1 vccd1 hold5025/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5036 _16934_/Q vssd1 vssd1 vccd1 vccd1 hold5036/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5047 _12157_/X vssd1 vssd1 vccd1 vccd1 _17209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4302 _10936_/X vssd1 vssd1 vccd1 vccd1 _16802_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4313 _17617_/Q vssd1 vssd1 vccd1 vccd1 hold4313/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput120 hold5876/X vssd1 vssd1 vccd1 vccd1 hold5877/A sky130_fd_sc_hd__buf_6
Xhold5058 _17637_/Q vssd1 vssd1 vccd1 vccd1 hold5058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4324 _09748_/X vssd1 vssd1 vccd1 vccd1 _16406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput131 hold5857/X vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_12
Xhold5069 _12256_/X vssd1 vssd1 vccd1 vccd1 _17242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput142 _13030_/A vssd1 vssd1 vccd1 vccd1 load_status[2] sky130_fd_sc_hd__buf_12
Xhold4335 _17183_/Q vssd1 vssd1 vccd1 vccd1 hold4335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4346 _13642_/X vssd1 vssd1 vccd1 vccd1 _17667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3601 _16734_/Q vssd1 vssd1 vccd1 vccd1 hold3601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3612 _11143_/Y vssd1 vssd1 vccd1 vccd1 _16871_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4357 _16408_/Q vssd1 vssd1 vccd1 vccd1 hold4357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3623 _13815_/Y vssd1 vssd1 vccd1 vccd1 _13816_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4368 _11437_/X vssd1 vssd1 vccd1 vccd1 _16969_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3634 _10581_/Y vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4379 _17125_/Q vssd1 vssd1 vccd1 vccd1 hold4379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3645 _16913_/Q vssd1 vssd1 vccd1 vccd1 hold3645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2900 _14253_/X vssd1 vssd1 vccd1 vccd1 _17927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2911 _18165_/Q vssd1 vssd1 vccd1 vccd1 hold2911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3656 _10036_/Y vssd1 vssd1 vccd1 vccd1 _16502_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2922 _14444_/X vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3667 _11161_/Y vssd1 vssd1 vccd1 vccd1 _16877_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3678 _16533_/Q vssd1 vssd1 vccd1 vccd1 hold3678/X sky130_fd_sc_hd__buf_1
Xhold2933 _15082_/X vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3689 _13822_/Y vssd1 vssd1 vccd1 vccd1 _17727_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 _15190_/X vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2955 _18136_/Q vssd1 vssd1 vccd1 vccd1 hold2955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2966 _15136_/X vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07957_ hold2764/X _07991_/A2 _07956_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07957_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2977 _17923_/Q vssd1 vssd1 vccd1 vccd1 hold2977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2988 _08180_/X vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2999 _18086_/Q vssd1 vssd1 vccd1 vccd1 hold2999/X sky130_fd_sc_hd__dlygate4sd3_1
X_07888_ hold756/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07888_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _09918_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09558_ _10098_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09558_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _15513_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09489_ _13048_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_109_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11520_ _12018_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _11640_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__or2_1
XFILLER_0_190_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10402_ hold4213/X _10646_/B _10401_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10402_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14170_ _15515_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14170_/X sky130_fd_sc_hd__or2_1
X_11382_ _11670_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__or2_1
X_13121_ _13121_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__and2_1
XFILLER_0_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10333_ hold4561/X _10619_/B _10332_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _10333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5570 _16843_/Q vssd1 vssd1 vccd1 vccd1 hold5570/X sky130_fd_sc_hd__dlygate4sd3_1
X_13052_ _17522_/Q _13056_/C _13056_/D _17523_/Q vssd1 vssd1 vccd1 vccd1 _13052_/X
+ sky130_fd_sc_hd__and4bb_4
X_10264_ hold4840/X _10589_/B _10263_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10264_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5581 _11371_/X vssd1 vssd1 vccd1 vccd1 _16947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5592 _16359_/Q vssd1 vssd1 vccd1 vccd1 hold5592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12003_ _13716_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4880 _11446_/X vssd1 vssd1 vccd1 vccd1 _16972_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10195_ hold5114/X _10073_/B _10194_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _10195_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4891 _16558_/Q vssd1 vssd1 vccd1 vccd1 hold4891/X sky130_fd_sc_hd__dlygate4sd3_1
X_17860_ _17862_/CLK hold984/X vssd1 vssd1 vccd1 vccd1 hold983/A sky130_fd_sc_hd__dfxtp_1
X_16811_ _18046_/CLK _16811_/D vssd1 vssd1 vccd1 vccd1 _16811_/Q sky130_fd_sc_hd__dfxtp_1
X_17791_ _17887_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout380 _14864_/B vssd1 vssd1 vccd1 vccd1 _14894_/B sky130_fd_sc_hd__buf_6
XFILLER_0_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout391 _14680_/Y vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__buf_6
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _15515_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13954_/X sky130_fd_sc_hd__or2_1
X_16742_ _18043_/CLK _16742_/D vssd1 vssd1 vccd1 vccd1 _16742_/Q sky130_fd_sc_hd__dfxtp_1
X_12905_ hold3201/X _12904_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12906_/B sky130_fd_sc_hd__mux2_1
X_16673_ _18231_/CLK _16673_/D vssd1 vssd1 vccd1 vccd1 _16673_/Q sky130_fd_sc_hd__dfxtp_1
X_13885_ _13888_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _13885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18412_ _18423_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ hold2340/X _12835_/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__mux2_1
X_15624_ _17844_/CLK _15624_/D vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18343_ _18416_/CLK hold431/X vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ hold800/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__or2_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12767_ hold3547/X _12766_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__mux2_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ hold1563/X _14554_/A2 _14505_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _14506_/X
+ sky130_fd_sc_hd__o211a_1
X_11718_ hold3182/X _12204_/A _11717_/X vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18274_ _18371_/CLK hold492/X vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_15486_ hold726/X _15486_/A2 _15486_/B1 hold673/X vssd1 vssd1 vccd1 vccd1 _15486_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ hold3412/X _12697_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17225_ _17257_/CLK _17225_/D vssd1 vssd1 vccd1 vccd1 _17225_/Q sky130_fd_sc_hd__dfxtp_1
X_14437_ _15551_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__or2_1
Xinput11 input11/A vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11649_/X sky130_fd_sc_hd__or2_1
Xinput22 input22/A vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 input33/A vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput44 input44/A vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
X_17156_ _17844_/CLK _17156_/D vssd1 vssd1 vccd1 vccd1 _17156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput55 input55/A vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
X_14368_ _14368_/A _14368_/B vssd1 vssd1 vccd1 vccd1 _17983_/D sky130_fd_sc_hd__and2_1
XFILLER_0_13_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold806 hold806/A vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _18410_/CLK _16107_/D vssd1 vssd1 vccd1 vccd1 hold691/A sky130_fd_sc_hd__dfxtp_1
Xhold817 hold817/A vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ hold1786/X _17560_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__mux2_1
Xhold828 hold828/A vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 hold839/A vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17087_ _18032_/CLK _17087_/D vssd1 vssd1 vccd1 vccd1 _17087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14299_ hold1061/X _14333_/A2 _14298_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _14299_/X
+ sky130_fd_sc_hd__o211a_1
X_16038_ _17340_/CLK _16038_/D vssd1 vssd1 vccd1 vccd1 hold718/A sky130_fd_sc_hd__dfxtp_1
X_08860_ hold359/X hold695/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__mux2_1
Xhold2207 _15690_/Q vssd1 vssd1 vccd1 vccd1 hold2207/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_177_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18066_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2218 _18106_/Q vssd1 vssd1 vccd1 vccd1 hold2218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 _09159_/X vssd1 vssd1 vccd1 vccd1 _16192_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07811_ hold925/X hold792/X hold898/X hold1771/X vssd1 vssd1 vccd1 vccd1 _07811_/X
+ sky130_fd_sc_hd__or4b_2
Xhold1506 _14617_/X vssd1 vssd1 vccd1 vccd1 _18102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18411_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1517 _17919_/Q vssd1 vssd1 vccd1 vccd1 hold1517/X sky130_fd_sc_hd__dlygate4sd3_1
X_08791_ hold14/X hold227/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__mux2_1
Xhold1528 _14945_/X vssd1 vssd1 vccd1 vccd1 _18259_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ _18060_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 hold422/A sky130_fd_sc_hd__dfxtp_1
Xhold1539 _14725_/X vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ _09438_/B _16292_/Q vssd1 vssd1 vccd1 vccd1 _09412_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09343_ hold784/X _15231_/A hold270/X hold241/X vssd1 vssd1 vccd1 vccd1 _09352_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _12756_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _16248_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _15559_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08225_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ hold624/A hold279/X hold606/X hold298/X vssd1 vssd1 vccd1 vccd1 _15492_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ hold837/X _08088_/B _08086_/Y _13939_/A vssd1 vssd1 vccd1 vccd1 hold838/A
+ sky130_fd_sc_hd__o211a_1
Xhold4110 _10312_/X vssd1 vssd1 vccd1 vccd1 _16594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4121 _17045_/Q vssd1 vssd1 vccd1 vccd1 hold4121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4132 _10687_/X vssd1 vssd1 vccd1 vccd1 _16719_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4143 _16588_/Q vssd1 vssd1 vccd1 vccd1 hold4143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4154 _11416_/X vssd1 vssd1 vccd1 vccd1 _16962_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4165 _16564_/Q vssd1 vssd1 vccd1 vccd1 hold4165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3420 _17140_/Q vssd1 vssd1 vccd1 vccd1 hold3420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3431 _16517_/Q vssd1 vssd1 vccd1 vccd1 hold3431/X sky130_fd_sc_hd__clkbuf_2
Xhold4176 _16883_/Q vssd1 vssd1 vccd1 vccd1 hold4176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3442 _16996_/Q vssd1 vssd1 vccd1 vccd1 hold3442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4187 _10915_/X vssd1 vssd1 vccd1 vccd1 _16795_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3453 _16617_/Q vssd1 vssd1 vccd1 vccd1 hold3453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4198 _16504_/Q vssd1 vssd1 vccd1 vccd1 hold4198/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3464 _09877_/X vssd1 vssd1 vccd1 vccd1 _16449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2730 _18173_/Q vssd1 vssd1 vccd1 vccd1 hold2730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3475 _11929_/X vssd1 vssd1 vccd1 vccd1 _17133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2741 _14317_/X vssd1 vssd1 vccd1 vccd1 _17958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3486 _17419_/Q vssd1 vssd1 vccd1 vccd1 hold3486/X sky130_fd_sc_hd__dlygate4sd3_1
X_08989_ hold44/X hold350/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08990_/B sky130_fd_sc_hd__mux2_1
Xhold3497 _17415_/Q vssd1 vssd1 vccd1 vccd1 hold3497/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2752 _16157_/Q vssd1 vssd1 vccd1 vccd1 hold2752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2763 _14169_/X vssd1 vssd1 vccd1 vccd1 _17887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2774 _18193_/Q vssd1 vssd1 vccd1 vccd1 hold2774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2785 _18081_/Q vssd1 vssd1 vccd1 vccd1 hold2785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2796 _08463_/X vssd1 vssd1 vccd1 vccd1 _15860_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ hold4039/X _11150_/B _10950_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10951_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13670_ hold2534/X _17677_/Q _13862_/C vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10882_ hold3232/X _11171_/B _10881_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10882_/X
+ sky130_fd_sc_hd__o211a_1
X_12621_ _12855_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _17383_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ hold645/X _15486_/A2 _15446_/B1 hold311/X vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__a22o_1
X_12552_ _12924_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _17360_/D sky130_fd_sc_hd__and2_1
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ hold4504/X _11798_/B _11502_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11503_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15271_ _16291_/Q _15477_/A2 _15487_/B1 hold496/X _15270_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/D sky130_fd_sc_hd__a221o_1
X_12483_ hold219/X _12509_/A2 _12505_/A3 _12482_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold220/A sky130_fd_sc_hd__o311a_1
X_17010_ _17889_/CLK _17010_/D vssd1 vssd1 vccd1 vccd1 _17010_/Q sky130_fd_sc_hd__dfxtp_1
X_14222_ _14972_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11434_ hold4834/X _11617_/A2 _11433_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ hold1627/X _14148_/B _14152_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11365_ hold4137/X _11747_/B _11364_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11365_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13104_ _13097_/X _13103_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17531_/D sky130_fd_sc_hd__o21a_1
X_10316_ hold1538/X hold4321/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__mux2_1
X_14084_ _15537_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14084_/X sky130_fd_sc_hd__or2_1
X_11296_ hold5560/X _11783_/B _11295_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11296_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _17523_/Q _13034_/X _13048_/A _13035_/D vssd1 vssd1 vccd1 vccd1 _13035_/X
+ sky130_fd_sc_hd__and4bb_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _18072_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_1
X_10247_ hold2141/X _16573_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_270_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17897_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17843_ _17873_/CLK hold774/X vssd1 vssd1 vccd1 vccd1 hold773/A sky130_fd_sc_hd__dfxtp_1
X_10178_ hold1732/X _16550_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__mux2_1
X_17774_ _17870_/CLK _17774_/D vssd1 vssd1 vccd1 vccd1 hold351/A sky130_fd_sc_hd__dfxtp_1
X_14986_ _14986_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ _18190_/CLK _16725_/D vssd1 vssd1 vccd1 vccd1 _16725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ _14350_/A _13937_/B vssd1 vssd1 vccd1 vccd1 _17776_/D sky130_fd_sc_hd__and2_1
X_16656_ _18214_/CLK _16656_/D vssd1 vssd1 vccd1 vccd1 _16656_/Q sky130_fd_sc_hd__dfxtp_1
X_13868_ _17743_/Q _13868_/B _13868_/C vssd1 vssd1 vccd1 vccd1 _13868_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12819_ _12825_/A _12819_/B vssd1 vssd1 vccd1 vccd1 _17449_/D sky130_fd_sc_hd__and2_1
X_15607_ _17453_/CLK _15607_/D vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16587_ _18268_/CLK _16587_/D vssd1 vssd1 vccd1 vccd1 _16587_/Q sky130_fd_sc_hd__dfxtp_1
X_13799_ hold1990/X hold3255/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__mux2_1
X_18326_ _18390_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ hold2367/X _15547_/B _15537_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _15538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15469_ _17322_/Q _15479_/A2 _09392_/B _16099_/Q _15468_/X vssd1 vssd1 vccd1 vccd1
+ _15471_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18257_ _18319_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ hold1278/X _08029_/B _08009_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _08010_/X
+ sky130_fd_sc_hd__o211a_1
X_17208_ _17208_/CLK _17208_/D vssd1 vssd1 vccd1 vccd1 _17208_/Q sky130_fd_sc_hd__dfxtp_1
X_18188_ _18220_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold603 la_data_in[28] vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold614 hold614/A vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17139_ _17865_/CLK _17139_/D vssd1 vssd1 vccd1 vccd1 _17139_/Q sky130_fd_sc_hd__dfxtp_1
Xhold625 hold625/A vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold636 hold664/X vssd1 vssd1 vccd1 vccd1 hold665/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 hold647/A vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _10055_/A _10601_/B _09960_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09961_/X
+ sky130_fd_sc_hd__o211a_1
Xhold669 hold669/A vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ hold8/X hold277/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08913_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_176_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _17817_/Q vssd1 vssd1 vccd1 vccd1 hold2004/X sky130_fd_sc_hd__dlygate4sd3_1
X_09892_ hold5512/X _10780_/A2 _09891_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _09892_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 _08016_/X vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2026 _17806_/Q vssd1 vssd1 vccd1 vccd1 hold2026/X sky130_fd_sc_hd__dlygate4sd3_1
X_08843_ _15473_/A _08843_/B vssd1 vssd1 vccd1 vccd1 _16040_/D sky130_fd_sc_hd__and2_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _14446_/X vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _08514_/X vssd1 vssd1 vccd1 vccd1 _15884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2048 _16166_/Q vssd1 vssd1 vccd1 vccd1 hold2048/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 _15116_/X vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _15518_/X vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 _14849_/X vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1336 _08239_/X vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _15482_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _16007_/D sky130_fd_sc_hd__and2_1
Xhold1347 _15532_/X vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 _14003_/X vssd1 vssd1 vccd1 vccd1 _17807_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 _15017_/X vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17292_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ hold2030/X _09325_/B _09325_/Y _14360_/A vssd1 vssd1 vccd1 vccd1 _09326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09257_ _15533_/A hold2378/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ hold2131/X _08213_/B _08207_/Y _08381_/A vssd1 vssd1 vccd1 vccd1 _08208_/X
+ sky130_fd_sc_hd__o211a_1
X_09188_ _15517_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _08139_/A hold370/X vssd1 vssd1 vccd1 vccd1 _15708_/D sky130_fd_sc_hd__and2_1
X_11150_ _16874_/Q _11150_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ _10485_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2_1
X_11081_ hold2828/X hold4159/X _11177_/C vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__mux2_1
Xhold3250 _11815_/X vssd1 vssd1 vccd1 vccd1 _17095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3261 _16631_/Q vssd1 vssd1 vccd1 vccd1 hold3261/X sky130_fd_sc_hd__dlygate4sd3_1
X_10032_ _13198_/A _09954_/A _10031_/X vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__a21oi_1
Xhold3272 _10447_/X vssd1 vssd1 vccd1 vccd1 _16639_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3283 _16405_/Q vssd1 vssd1 vccd1 vccd1 hold3283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3294 _13339_/X vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2560 _14915_/X vssd1 vssd1 vccd1 vccd1 _18244_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14840_ _15233_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__or2_1
Xhold2571 _14891_/X vssd1 vssd1 vccd1 vccd1 _18234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2582 _16163_/Q vssd1 vssd1 vccd1 vccd1 hold2582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2593 _14621_/X vssd1 vssd1 vccd1 vccd1 _18104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1870 _17940_/Q vssd1 vssd1 vccd1 vccd1 hold1870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1881 _17850_/Q vssd1 vssd1 vccd1 vccd1 hold1881/X sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ hold2668/X _14774_/B _14770_/Y _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14771_/X
+ sky130_fd_sc_hd__o211a_1
X_11983_ hold4335/X _13844_/B _11982_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _11983_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1892 _08196_/X vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13722_ _13800_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13722_/X sky130_fd_sc_hd__or2_1
X_16510_ _18385_/CLK _16510_/D vssd1 vssd1 vccd1 vccd1 _16510_/Q sky130_fd_sc_hd__dfxtp_1
X_10934_ hold2491/X _16802_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__mux2_1
X_17490_ _17517_/CLK _17490_/D vssd1 vssd1 vccd1 vccd1 _17490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ _18386_/CLK _16441_/D vssd1 vssd1 vccd1 vccd1 _16441_/Q sky130_fd_sc_hd__dfxtp_1
X_13653_ _13779_/A _13653_/B vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ hold2490/X _16779_/Q _11066_/S vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ hold2594/X hold3253/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__mux2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _18363_/CLK _16372_/D vssd1 vssd1 vccd1 vccd1 _16372_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13770_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10796_ hold1553/X hold4771/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__mux2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15490_/A1 _15315_/X _15322_/X _15490_/B1 hold5843/A vssd1 vssd1 vccd1 vccd1
+ _15323_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _18267_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ hold1067/X hold3586/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15254_ _15414_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__and2_1
X_18042_ _18042_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ _17326_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ hold843/X _14202_/B _14204_/X _13939_/A vssd1 vssd1 vccd1 vccd1 hold844/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ hold993/X _16963_/Q _12341_/C vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15185_ _15185_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__or2_1
X_12397_ hold126/X hold457/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ _14529_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14136_/X sky130_fd_sc_hd__or2_1
X_11348_ hold1235/X _16940_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ hold2503/X _14105_/A2 _14066_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _14067_/X
+ sky130_fd_sc_hd__o211a_1
X_11279_ _17765_/Q hold5365/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__mux2_1
X_13018_ hold1868/X _13003_/Y _13017_/X _12936_/A vssd1 vssd1 vccd1 vccd1 _13018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _17889_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _18073_/CLK _17757_/D vssd1 vssd1 vccd1 vccd1 _17757_/Q sky130_fd_sc_hd__dfxtp_1
X_14969_ hold2618/X _15006_/B _14968_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _14969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16708_ _18071_/CLK _16708_/D vssd1 vssd1 vccd1 vccd1 _16708_/Q sky130_fd_sc_hd__dfxtp_1
X_08490_ hold730/X _08498_/B vssd1 vssd1 vccd1 vccd1 _08490_/X sky130_fd_sc_hd__or2_1
X_17688_ _17725_/CLK _17688_/D vssd1 vssd1 vccd1 vccd1 _17688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _18131_/CLK _16639_/D vssd1 vssd1 vccd1 vccd1 _16639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ hold1507/X _09119_/A2 _09110_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09111_/X
+ sky130_fd_sc_hd__o211a_1
X_18309_ _18334_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09042_ hold8/X hold512/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_192_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18055_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold411 hold411/A vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold422/A vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 hold444/A vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold455 hold455/A vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__clkbuf_8
Xhold477 hold477/A vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 hold784/X vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__buf_8
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09944_ hold2748/X hold3285/X _10571_/C vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__mux2_1
Xhold499 input9/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 hold770/X vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__buf_8
XFILLER_0_99_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout924 hold891/X vssd1 vssd1 vccd1 vccd1 _14970_/A sky130_fd_sc_hd__buf_4
Xfanout935 hold1452/X vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__buf_4
Xfanout946 hold943/X vssd1 vssd1 vccd1 vccd1 hold944/A sky130_fd_sc_hd__buf_6
X_09875_ hold1063/X _16449_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _08420_/X vssd1 vssd1 vccd1 vccd1 _15840_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _14821_/X vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ hold136/X hold165/X _08860_/S vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__mux2_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _17805_/Q vssd1 vssd1 vccd1 vccd1 hold1122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _14045_/X vssd1 vssd1 vccd1 vccd1 _17828_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _17922_/Q vssd1 vssd1 vccd1 vccd1 hold1144/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _14438_/X vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 _13971_/X vssd1 vssd1 vccd1 vccd1 _17792_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ hold59/X hold706/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__mux2_1
Xhold1177 _15761_/Q vssd1 vssd1 vccd1 vccd1 hold1177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _08410_/X vssd1 vssd1 vccd1 vccd1 _15835_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _18037_/Q vssd1 vssd1 vccd1 vccd1 hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _15244_/A hold427/X vssd1 vssd1 vccd1 vccd1 _15965_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ hold3126/X _10554_/A _10649_/X vssd1 vssd1 vccd1 vccd1 _10650_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09309_ _15531_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ hold3633/X _10485_/A _10580_/X vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _17264_/Q _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_209_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17896_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12251_ hold2687/X _17241_/Q _13388_/S vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11202_ hold5309/X _11106_/A _11201_/X vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ hold1359/X hold4737/X _13844_/C vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__mux2_1
X_11133_ _11640_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16990_ _17870_/CLK _16990_/D vssd1 vssd1 vccd1 vccd1 _16990_/Q sky130_fd_sc_hd__dfxtp_1
X_15941_ _17292_/CLK _15941_/D vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__dfxtp_1
X_11064_ _11067_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__or2_1
Xhold3080 _17457_/Q vssd1 vssd1 vccd1 vccd1 hold3080/X sky130_fd_sc_hd__dlygate4sd3_1
X_10015_ _11203_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10015_/Y sky130_fd_sc_hd__nor2_1
Xhold3091 _17454_/Q vssd1 vssd1 vccd1 vccd1 hold3091/X sky130_fd_sc_hd__dlygate4sd3_1
X_15872_ _17583_/CLK hold876/X vssd1 vssd1 vccd1 vccd1 hold875/A sky130_fd_sc_hd__dfxtp_1
Xhold2390 _18348_/Q vssd1 vssd1 vccd1 vccd1 hold2390/X sky130_fd_sc_hd__dlygate4sd3_1
X_17611_ _17734_/CLK _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
X_14823_ hold2022/X _14822_/B _14822_/Y _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14823_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _18358_/CLK _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14754_ _14986_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14754_/X sky130_fd_sc_hd__or2_1
X_11966_ hold1455/X hold4846/X _13388_/S vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13705_ hold3255/X _13808_/B _13704_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13705_/X
+ sky130_fd_sc_hd__o211a_1
X_10917_ _11115_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__or2_1
X_14685_ hold1515/X _14720_/B _14684_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14685_/X
+ sky130_fd_sc_hd__o211a_1
X_17473_ _17475_/CLK _17473_/D vssd1 vssd1 vccd1 vccd1 _17473_/Q sky130_fd_sc_hd__dfxtp_1
X_11897_ hold2611/X hold3767/X _12377_/C vssd1 vssd1 vccd1 vccd1 _11898_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13636_ hold4238/X _13829_/B _13635_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13636_/X
+ sky130_fd_sc_hd__o211a_1
X_16424_ _18337_/CLK _16424_/D vssd1 vssd1 vccd1 vccd1 _16424_/Q sky130_fd_sc_hd__dfxtp_1
X_10848_ _11136_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16355_ _18388_/CLK _16355_/D vssd1 vssd1 vccd1 vccd1 _16355_/Q sky130_fd_sc_hd__dfxtp_1
X_13567_ hold5201/X _13883_/B _13566_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15306_ _17334_/Q _09362_/C _09362_/D hold459/X vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__a22o_1
X_12518_ hold3415/X _12517_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16286_ _18461_/CLK _16286_/D vssd1 vssd1 vccd1 vccd1 _16286_/Q sky130_fd_sc_hd__dfxtp_1
X_13498_ hold5110/X _13880_/B _13497_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13498_/X
+ sky130_fd_sc_hd__o211a_1
X_18025_ _18025_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
X_12449_ hold68/X _12509_/A2 _12505_/A3 _12448_/X _12420_/A vssd1 vssd1 vccd1 vccd1
+ hold69/A sky130_fd_sc_hd__o311a_1
X_15237_ _16132_/Q _09357_/A _15484_/B1 hold191/X _15236_/X vssd1 vssd1 vccd1 vccd1
+ _15242_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_23_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4709 _13750_/X vssd1 vssd1 vccd1 vccd1 _17703_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15168_ hold1962/X hold609/X _15167_/Y _15168_/C1 vssd1 vssd1 vccd1 vccd1 _15168_/X
+ sky130_fd_sc_hd__o211a_1
X_14119_ hold1077/X hold587/X _14118_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14119_/X
+ sky130_fd_sc_hd__o211a_1
X_15099_ _15099_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15099_/X sky130_fd_sc_hd__or2_1
X_07990_ _14786_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__or2_1
Xfanout209 _09494_/X vssd1 vssd1 vccd1 vccd1 fanout209/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09660_ _09954_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08611_ hold26/X hold368/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__mux2_1
X_17809_ _17873_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_1
X_09591_ _09975_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__or2_1
X_08542_ hold41/X hold533/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08473_ hold1397/X _08486_/B _08472_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _08473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_302_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17694_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_190_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09025_ _15491_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _16129_/D sky130_fd_sc_hd__and2_1
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5900 _16528_/Q vssd1 vssd1 vccd1 vccd1 hold5900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5911 _17546_/Q vssd1 vssd1 vccd1 vccd1 hold5911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5922 _17551_/Q vssd1 vssd1 vccd1 vccd1 hold5922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5933 _17534_/Q vssd1 vssd1 vccd1 vccd1 hold5933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5944 hold6007/X vssd1 vssd1 vccd1 vccd1 hold5944/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold230 input31/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5955 _15672_/Q vssd1 vssd1 vccd1 vccd1 hold5955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold654/X vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__clkbuf_4
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5966 _18073_/Q vssd1 vssd1 vccd1 vccd1 hold5966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5977 _18433_/Q vssd1 vssd1 vccd1 vccd1 hold5977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5988 data_in[19] vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 input44/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5999 _18419_/Q vssd1 vssd1 vccd1 vccd1 hold5999/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__clkbuf_2
Xhold285 input5/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 input58/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _08970_/A vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__clkbuf_4
Xfanout721 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__buf_4
Xfanout732 _15364_/A vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__clkbuf_4
X_09927_ _09987_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout743 _08111_/A vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__buf_4
Xfanout754 _14378_/A vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__buf_4
Xfanout765 _13753_/C1 vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__buf_4
Xfanout776 _12274_/C1 vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__buf_4
X_09858_ _09954_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__or2_1
Xfanout787 _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__buf_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 _15072_/A vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__buf_4
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _09011_/A hold661/X vssd1 vssd1 vccd1 vccd1 _16023_/D sky130_fd_sc_hd__and2_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09789_ _09987_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__or2_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ _12204_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _15103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_125 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ hold5281/X _12234_/A _11750_/X vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ hold4771/X _11192_/B _10701_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10702_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ hold820/X _14481_/B _14469_/X _13935_/A vssd1 vssd1 vccd1 vccd1 hold821/A
+ sky130_fd_sc_hd__o211a_1
X_11682_ _12036_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ hold1640/X _17594_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10633_ _10651_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _10633_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_165_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16140_ _17523_/CLK _16140_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ hold2795/X hold3690/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__mux2_1
X_10564_ hold3545/X _10568_/B _10563_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _16678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ hold3808/X _13716_/A _12302_/X vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__a21oi_1
X_16071_ _17318_/CLK _16071_/D vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__dfxtp_1
X_13283_ _13282_/X hold5889/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__mux2_1
X_10495_ hold4252/X _10589_/B _10494_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10495_/X
+ sky130_fd_sc_hd__o211a_1
X_15022_ _15030_/A _15022_/B vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__and2_1
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _12267_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ hold5464/X _11210_/B _11115_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _11116_/X
+ sky130_fd_sc_hd__o211a_1
X_12096_ _13797_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__or2_1
X_16973_ _17856_/CLK _16973_/D vssd1 vssd1 vccd1 vccd1 _16973_/Q sky130_fd_sc_hd__dfxtp_1
X_15924_ _18406_/CLK _15924_/D vssd1 vssd1 vccd1 vccd1 hold677/A sky130_fd_sc_hd__dfxtp_1
X_11047_ hold4026/X _11150_/B _11046_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _11047_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 input9/A vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _17686_/CLK _15855_/D vssd1 vssd1 vccd1 vccd1 _15855_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14984_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__or2_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _17745_/CLK hold817/X vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12998_ hold3456/X _12997_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__mux2_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _17525_/CLK _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ hold2793/X _14774_/B _14736_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14737_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ _12255_/A _11949_/B vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__or2_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17456_ _17456_/CLK _17456_/D vssd1 vssd1 vccd1 vccd1 _17456_/Q sky130_fd_sc_hd__dfxtp_1
X_14668_ _15169_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16407_ _18390_/CLK _16407_/D vssd1 vssd1 vccd1 vccd1 _16407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13619_ hold1877/X hold4557/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13620_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17387_ _18438_/CLK _17387_/D vssd1 vssd1 vccd1 vccd1 _17387_/Q sky130_fd_sc_hd__dfxtp_1
X_14599_ hold1809/X _14610_/B _14598_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _14599_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16338_ _18373_/CLK _16338_/D vssd1 vssd1 vccd1 vccd1 _16338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5207 _17684_/Q vssd1 vssd1 vccd1 vccd1 hold5207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5218 _15443_/X vssd1 vssd1 vccd1 vccd1 _15444_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16269_ _17981_/CLK _16269_/D vssd1 vssd1 vccd1 vccd1 _16269_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5229 _11758_/Y vssd1 vssd1 vccd1 vccd1 _17076_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18042_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4506 _16901_/Q vssd1 vssd1 vccd1 vccd1 hold4506/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4517 _10219_/X vssd1 vssd1 vccd1 vccd1 _16563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4528 _16407_/Q vssd1 vssd1 vccd1 vccd1 hold4528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4539 _11587_/X vssd1 vssd1 vccd1 vccd1 _17019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3805 _17104_/Q vssd1 vssd1 vccd1 vccd1 hold3805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3816 _13867_/Y vssd1 vssd1 vccd1 vccd1 _17742_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3827 _12319_/Y vssd1 vssd1 vccd1 vccd1 _17263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3838 _16351_/Q vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3849 _16724_/Q vssd1 vssd1 vccd1 vccd1 hold3849/X sky130_fd_sc_hd__dlygate4sd3_1
X_07973_ hold2044/X _07978_/B _07972_/Y _08171_/A vssd1 vssd1 vccd1 vccd1 _07973_/X
+ sky130_fd_sc_hd__o211a_1
X_09712_ hold5625/X _09992_/B _09711_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09712_/X
+ sky130_fd_sc_hd__o211a_1
X_09643_ hold5482/X _10025_/B _09642_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09643_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ hold4081/X _10571_/B _09573_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09574_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _15491_/A hold600/X vssd1 vssd1 vccd1 vccd1 _15887_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08456_ _14850_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08456_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _15825_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09008_ hold32/X hold372/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5730 _11479_/X vssd1 vssd1 vccd1 vccd1 _16983_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10280_ hold2907/X hold3487/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5741 _16847_/Q vssd1 vssd1 vccd1 vccd1 hold5741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5752 output94/X vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_12
Xhold5763 hold5910/X vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__buf_1
Xhold5774 output99/X vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_12
Xhold5785 hold5922/X vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold5796 output78/X vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_12
Xfanout540 _12445_/B vssd1 vssd1 vccd1 vccd1 _08999_/B sky130_fd_sc_hd__clkbuf_8
Xfanout551 hold121/X vssd1 vssd1 vccd1 vccd1 _08390_/S sky130_fd_sc_hd__clkbuf_8
Xfanout562 hold195/X vssd1 vssd1 vccd1 vccd1 _08152_/S sky130_fd_sc_hd__clkbuf_8
Xfanout573 _07924_/B vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__buf_6
X_13970_ _15531_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__or2_1
Xfanout584 _13057_/X vssd1 vssd1 vccd1 vccd1 _13306_/S sky130_fd_sc_hd__buf_8
Xfanout595 _12679_/S vssd1 vssd1 vccd1 vccd1 _12676_/S sky130_fd_sc_hd__buf_6
X_12921_ _12924_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _17483_/D sky130_fd_sc_hd__and2_1
X_15640_ _17205_/CLK _15640_/D vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12855_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _17460_/D sky130_fd_sc_hd__and2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ _12343_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11803_/Y sky130_fd_sc_hd__nor2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12789_/A _12783_/B vssd1 vssd1 vccd1 vccd1 _17437_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_295_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17275_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15571_ _17907_/CLK _15571_/D vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _18410_/CLK _17310_/D vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__dfxtp_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _12301_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11734_/Y sky130_fd_sc_hd__nor2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ hold2713/X _14541_/B _14521_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14522_/X
+ sky130_fd_sc_hd__o211a_1
X_18290_ _18358_/CLK hold776/X vssd1 vssd1 vccd1 vccd1 hold775/A sky130_fd_sc_hd__dfxtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_224_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17777_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17703_/CLK _17241_/D vssd1 vssd1 vccd1 vccd1 _17241_/Q sky130_fd_sc_hd__dfxtp_1
X_11665_ _11759_/A _12341_/B _11664_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11665_/X
+ sky130_fd_sc_hd__o211a_1
X_14453_ _14740_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ _13788_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10616_ _16696_/Q _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__and3_1
X_17172_ _17274_/CLK _17172_/D vssd1 vssd1 vccd1 vccd1 _17172_/Q sky130_fd_sc_hd__dfxtp_1
X_14384_ _14384_/A _14384_/B vssd1 vssd1 vccd1 vccd1 _17991_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11596_ hold4099/X _12329_/B _11595_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11596_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ _17531_/CLK _16123_/D vssd1 vssd1 vccd1 vccd1 hold374/A sky130_fd_sc_hd__dfxtp_1
X_13335_ _13800_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__or2_1
X_10547_ hold758/X hold4071/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16054_ _17307_/CLK _16054_/D vssd1 vssd1 vccd1 vccd1 _16054_/Q sky130_fd_sc_hd__dfxtp_1
X_13266_ _17584_/Q _17118_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13266_/X sky130_fd_sc_hd__mux2_1
X_10478_ hold2603/X _16650_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15005_ hold2524/X _15004_/B _15004_/Y _15070_/A vssd1 vssd1 vccd1 vccd1 _15005_/X
+ sky130_fd_sc_hd__o211a_1
X_12217_ hold4951/X _12311_/B _12216_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _12217_/X
+ sky130_fd_sc_hd__o211a_1
X_13197_ _13196_/X hold3678/X _13197_/S vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__mux2_1
X_12148_ hold5126/X _12362_/B _12147_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _12148_/X
+ sky130_fd_sc_hd__o211a_1
X_12079_ hold4482/X _13844_/B _12078_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12079_/X
+ sky130_fd_sc_hd__o211a_1
X_16956_ _17887_/CLK _16956_/D vssd1 vssd1 vccd1 vccd1 _16956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15907_ _17345_/CLK _15907_/D vssd1 vssd1 vccd1 vccd1 hold651/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16887_ _18067_/CLK _16887_/D vssd1 vssd1 vccd1 vccd1 _16887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _17697_/CLK _15838_/D vssd1 vssd1 vccd1 vccd1 _15838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15769_ _17725_/CLK _15769_/D vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08310_ hold2201/X _08323_/B _08309_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _08310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17508_ _17517_/CLK _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09290_ hold1471/X _09338_/A2 _09289_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08241_ hold2772/X _08262_/B _08240_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08241_/X
+ sky130_fd_sc_hd__o211a_1
X_17439_ _17439_/CLK _17439_/D vssd1 vssd1 vccd1 vccd1 _17439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_14 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _13260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _15519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ hold624/A hold279/X hold606/A hold298/A vssd1 vssd1 vccd1 vccd1 _15182_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA_58 _14866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 hold747/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5004 _11320_/X vssd1 vssd1 vccd1 vccd1 _16930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5015 _17195_/Q vssd1 vssd1 vccd1 vccd1 hold5015/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5026 _17167_/Q vssd1 vssd1 vccd1 vccd1 hold5026/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5037 _11236_/X vssd1 vssd1 vccd1 vccd1 _16902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5048 _16479_/Q vssd1 vssd1 vccd1 vccd1 hold5048/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput110 hold5835/X vssd1 vssd1 vccd1 vccd1 hold5836/A sky130_fd_sc_hd__buf_6
Xhold4303 _17066_/Q vssd1 vssd1 vccd1 vccd1 hold4303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4314 _13396_/X vssd1 vssd1 vccd1 vccd1 _17585_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput121 hold5858/X vssd1 vssd1 vccd1 vccd1 hold5859/A sky130_fd_sc_hd__buf_6
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5059 _13456_/X vssd1 vssd1 vccd1 vccd1 _17605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4325 _17696_/Q vssd1 vssd1 vccd1 vccd1 hold4325/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput132 hold4842/X vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput143 hold1551/X vssd1 vssd1 vccd1 vccd1 load_status[3] sky130_fd_sc_hd__buf_12
XFILLER_0_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4336 _11983_/X vssd1 vssd1 vccd1 vccd1 _17151_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17878_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4347 _17731_/Q vssd1 vssd1 vccd1 vccd1 hold4347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3602 _11211_/Y vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3613 _16925_/Q vssd1 vssd1 vccd1 vccd1 hold3613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4358 _09658_/X vssd1 vssd1 vccd1 vccd1 _16376_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3624 _13816_/Y vssd1 vssd1 vccd1 vccd1 _17725_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4369 _16941_/Q vssd1 vssd1 vccd1 vccd1 hold4369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3635 _10582_/Y vssd1 vssd1 vccd1 vccd1 _16684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2901 _18171_/Q vssd1 vssd1 vccd1 vccd1 hold2901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3646 _11748_/Y vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2912 _14749_/X vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3657 _16014_/Q vssd1 vssd1 vccd1 vccd1 _15445_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3668 hold5864/X vssd1 vssd1 vccd1 vccd1 hold5865/A sky130_fd_sc_hd__buf_4
Xhold2923 _18247_/Q vssd1 vssd1 vccd1 vccd1 hold2923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3679 _10608_/Y vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 _18435_/Q vssd1 vssd1 vccd1 vccd1 hold2934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2945 _16173_/Q vssd1 vssd1 vccd1 vccd1 hold2945/X sky130_fd_sc_hd__dlygate4sd3_1
X_07956_ _15525_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07956_/X sky130_fd_sc_hd__or2_1
Xhold2956 _14689_/X vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2967 _18046_/Q vssd1 vssd1 vccd1 vccd1 hold2967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2978 _14245_/X vssd1 vssd1 vccd1 vccd1 _17923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2989 _17751_/Q vssd1 vssd1 vccd1 vccd1 hold2989/X sky130_fd_sc_hd__dlygate4sd3_1
X_07887_ hold1284/X _07918_/B _07886_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _07887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ hold2487/X _16366_/Q _09893_/S vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__mux2_1
X_09557_ hold1659/X _13214_/A _10601_/C vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08508_ hold962/X _08503_/Y _08507_/X _08161_/A vssd1 vssd1 vccd1 vccd1 hold963/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _13046_/A _13035_/D vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08439_ _15553_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08439_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ hold1167/X hold4087/X _11735_/C vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10521_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__or2_1
X_11381_ hold2125/X hold5711/X _11765_/C vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13120_ _13113_/X _13119_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17533_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_15_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10332_ _10524_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ _13051_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and2_1
Xhold5560 _16954_/Q vssd1 vssd1 vccd1 vccd1 hold5560/X sky130_fd_sc_hd__dlygate4sd3_1
X_10263_ _10551_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__or2_1
Xhold5571 _10963_/X vssd1 vssd1 vccd1 vccd1 _16811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5582 _16670_/Q vssd1 vssd1 vccd1 vccd1 hold5582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5593 _09511_/X vssd1 vssd1 vccd1 vccd1 _16327_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12002_ hold1278/X _17158_/Q _13811_/C vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__mux2_1
Xhold4870 _12085_/X vssd1 vssd1 vccd1 vccd1 _17185_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10194_ _10506_/A _10194_/B vssd1 vssd1 vccd1 vccd1 _10194_/X sky130_fd_sc_hd__or2_1
Xhold4881 _17030_/Q vssd1 vssd1 vccd1 vccd1 hold4881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4892 _10108_/X vssd1 vssd1 vccd1 vccd1 _16526_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16810_ _18013_/CLK _16810_/D vssd1 vssd1 vccd1 vccd1 _16810_/Q sky130_fd_sc_hd__dfxtp_1
X_17790_ _18051_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout370 _15109_/B vssd1 vssd1 vccd1 vccd1 _15113_/B sky130_fd_sc_hd__buf_6
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout381 _14842_/Y vssd1 vssd1 vccd1 vccd1 _14882_/B sky130_fd_sc_hd__buf_8
X_16741_ _18042_/CLK _16741_/D vssd1 vssd1 vccd1 vccd1 _16741_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout392 _14668_/B vssd1 vssd1 vccd1 vccd1 _14678_/B sky130_fd_sc_hd__clkbuf_8
X_13953_ hold2895/X _13980_/B _13952_/X _12666_/A vssd1 vssd1 vccd1 vccd1 _13953_/X
+ sky130_fd_sc_hd__o211a_1
X_12904_ hold1840/X hold3001/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__mux2_1
X_16672_ _18230_/CLK _16672_/D vssd1 vssd1 vccd1 vccd1 _16672_/Q sky130_fd_sc_hd__dfxtp_1
X_13884_ hold4544/X _13788_/A _13883_/X vssd1 vssd1 vccd1 vccd1 _13884_/Y sky130_fd_sc_hd__a21oi_1
X_18411_ _18411_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
X_15623_ _17279_/CLK _15623_/D vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _16224_/Q _17456_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__mux2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18420_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ hold2437/X _15547_/B _15553_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _15554_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ hold2120/X hold3406/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14970_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _17063_/Q _12299_/B _11717_/C vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__and3_1
X_18273_ _18273_/CLK hold686/X vssd1 vssd1 vccd1 vccd1 hold685/A sky130_fd_sc_hd__dfxtp_1
X_15485_ hold694/X _15485_/A2 _15485_/B1 hold727/X vssd1 vssd1 vccd1 vccd1 _15485_/X
+ sky130_fd_sc_hd__a22o_1
X_12697_ hold3003/X hold3410/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
X_17224_ _17453_/CLK _17224_/D vssd1 vssd1 vccd1 vccd1 _17224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ hold1661/X _17040_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__mux2_1
X_14436_ hold2052/X _14433_/B _14435_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _14436_/X
+ sky130_fd_sc_hd__o211a_1
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
Xinput23 input23/A vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 input34/A vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 input45/A vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_17155_ _17283_/CLK _17155_/D vssd1 vssd1 vccd1 vccd1 _17155_/Q sky130_fd_sc_hd__dfxtp_1
X_11579_ hold2551/X hold3890/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11580_/B sky130_fd_sc_hd__mux2_1
X_14367_ _15535_/A hold1722/X hold275/X vssd1 vssd1 vccd1 vccd1 _14368_/B sky130_fd_sc_hd__mux2_1
Xinput56 input56/A vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xhold807 hold807/A vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 input67/A vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _18417_/CLK _16106_/D vssd1 vssd1 vccd1 vccd1 _16106_/Q sky130_fd_sc_hd__dfxtp_1
Xhold818 hold818/A vssd1 vssd1 vccd1 vccd1 hold818/X sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ hold3313/X _13814_/B _13317_/X _13627_/C1 vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__o211a_1
X_17086_ _17870_/CLK _17086_/D vssd1 vssd1 vccd1 vccd1 _17086_/Q sky130_fd_sc_hd__dfxtp_1
Xhold829 hold829/A vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ hold826/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16037_ _17513_/CLK _16037_/D vssd1 vssd1 vccd1 vccd1 hold420/A sky130_fd_sc_hd__dfxtp_1
X_13249_ _13249_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__and2_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2208 _08101_/X vssd1 vssd1 vccd1 vccd1 _15690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2219 _14625_/X vssd1 vssd1 vccd1 vccd1 _18106_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07810_ _12442_/A _17751_/Q vssd1 vssd1 vccd1 vccd1 _07810_/Y sky130_fd_sc_hd__nand2_1
X_08790_ _15482_/A hold381/X vssd1 vssd1 vccd1 vccd1 _16015_/D sky130_fd_sc_hd__and2_1
Xhold1507 _16170_/Q vssd1 vssd1 vccd1 vccd1 hold1507/X sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ _18020_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 hold483/A sky130_fd_sc_hd__dfxtp_1
Xhold1518 _14237_/X vssd1 vssd1 vccd1 vccd1 _17919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _18436_/Q vssd1 vssd1 vccd1 vccd1 hold1529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16939_ _17852_/CLK _16939_/D vssd1 vssd1 vccd1 vccd1 _16939_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_146_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09411_ _07785_/Y _09447_/A _15314_/A _09410_/X vssd1 vssd1 vccd1 vccd1 _09411_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ _15549_/A hold1863/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ hold2814/X _08209_/B _08223_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08155_ _15498_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08086_ _14950_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4100 _11596_/X vssd1 vssd1 vccd1 vccd1 _17022_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4111 _16374_/Q vssd1 vssd1 vccd1 vccd1 hold4111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4122 _11569_/X vssd1 vssd1 vccd1 vccd1 _17013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4133 _17082_/Q vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4144 _10198_/X vssd1 vssd1 vccd1 vccd1 _16556_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4155 _16620_/Q vssd1 vssd1 vccd1 vccd1 hold4155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3410 _17410_/Q vssd1 vssd1 vccd1 vccd1 hold3410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4166 _10126_/X vssd1 vssd1 vccd1 vccd1 _16532_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3421 _11854_/X vssd1 vssd1 vccd1 vccd1 _17108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3432 _10561_/X vssd1 vssd1 vccd1 vccd1 _16677_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4177 _11083_/X vssd1 vssd1 vccd1 vccd1 _16851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4188 _16591_/Q vssd1 vssd1 vccd1 vccd1 hold4188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3443 _11422_/X vssd1 vssd1 vccd1 vccd1 _16964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3454 _10285_/X vssd1 vssd1 vccd1 vccd1 _16585_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4199 _09946_/X vssd1 vssd1 vccd1 vccd1 _16472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2720 _14985_/X vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3465 _17351_/Q vssd1 vssd1 vccd1 vccd1 hold3465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2731 _14765_/X vssd1 vssd1 vccd1 vccd1 _18173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3476 _17429_/Q vssd1 vssd1 vccd1 vccd1 hold3476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3487 _16584_/Q vssd1 vssd1 vccd1 vccd1 hold3487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2742 _17930_/Q vssd1 vssd1 vccd1 vccd1 hold2742/X sky130_fd_sc_hd__dlygate4sd3_1
X_08988_ _09003_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _16111_/D sky130_fd_sc_hd__and2_1
Xhold3498 _17691_/Q vssd1 vssd1 vccd1 vccd1 hold3498/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2753 _09085_/X vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2764 _15621_/Q vssd1 vssd1 vccd1 vccd1 hold2764/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2775 _14807_/X vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2786 _14575_/X vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07939_ _14735_/A _08504_/A vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__or2_4
Xhold2797 _18161_/Q vssd1 vssd1 vccd1 vccd1 hold2797/X sky130_fd_sc_hd__dlygate4sd3_1
X_10950_ _11061_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/X sky130_fd_sc_hd__or2_1
X_09609_ _11067_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__or2_1
X_10881_ _11076_/A _10881_/B vssd1 vssd1 vccd1 vccd1 _10881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ hold3020/X _12619_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ hold3297/X _12550_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _12153_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15270_ hold719/X _09367_/A _09392_/A hold593/X vssd1 vssd1 vccd1 vccd1 _15270_/X
+ sky130_fd_sc_hd__a22o_1
X_12482_ _17334_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11433_ _11616_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__or2_1
X_14221_ hold1652/X _14216_/Y _14220_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _14221_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14152_ _15551_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11364_ _11652_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ hold4435/X _10619_/B _10314_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _10315_/X
+ sky130_fd_sc_hd__o211a_1
X_13103_ _13183_/A1 _13101_/X _13102_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__o211a_1
X_14083_ hold1686/X _14094_/B _14082_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__o211a_1
X_11295_ _12051_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__or2_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13053_/A _13056_/C _17520_/Q _13034_/D vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__and4_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _18072_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5390 _11101_/X vssd1 vssd1 vccd1 vccd1 _16857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10246_ hold3326/X _10610_/B _10245_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10246_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17842_ _17905_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_1
X_10177_ hold4858/X _10571_/B _10176_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _10177_/X
+ sky130_fd_sc_hd__o211a_1
X_17773_ _17901_/CLK _17773_/D vssd1 vssd1 vccd1 vccd1 hold402/A sky130_fd_sc_hd__dfxtp_1
X_14985_ hold2719/X _15004_/B _14984_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _14985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16724_ _18055_/CLK _16724_/D vssd1 vssd1 vccd1 vccd1 _16724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13936_ _14330_/A hold1334/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13937_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_159_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16655_ _18192_/CLK _16655_/D vssd1 vssd1 vccd1 vccd1 _16655_/Q sky130_fd_sc_hd__dfxtp_1
X_13867_ _13873_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _13867_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _17592_/CLK _15606_/D vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ hold3506/X _12817_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12819_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16586_ _18176_/CLK _16586_/D vssd1 vssd1 vccd1 vccd1 _16586_/Q sky130_fd_sc_hd__dfxtp_1
X_13798_ hold4256/X _12308_/B _13797_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _17719_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18325_ _18389_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _15537_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__or2_1
X_12749_ hold3027/X _12748_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18256_ _18360_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15468_ hold601/X _09367_/A _15486_/B1 hold660/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _17216_/CLK _17207_/D vssd1 vssd1 vccd1 vccd1 _17207_/Q sky130_fd_sc_hd__dfxtp_1
X_14419_ _15099_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ _18233_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15399_ hold312/X _09365_/B _15447_/B1 hold167/X _15398_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 hold604/A vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
X_17138_ _17170_/CLK _17138_/D vssd1 vssd1 vccd1 vccd1 _17138_/Q sky130_fd_sc_hd__dfxtp_1
Xhold615 hold626/X vssd1 vssd1 vccd1 vccd1 hold627/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 slv_done vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 hold666/X vssd1 vssd1 vccd1 vccd1 hold667/A sky130_fd_sc_hd__buf_6
Xhold648 hold648/A vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _10098_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__or2_1
Xhold659 hold659/A vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _18073_/CLK _17069_/D vssd1 vssd1 vccd1 vccd1 _17069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _12422_/A hold260/X vssd1 vssd1 vccd1 vccd1 _16073_/D sky130_fd_sc_hd__and2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _10779_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__or2_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _14023_/X vssd1 vssd1 vccd1 vccd1 _17817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2016 _18233_/Q vssd1 vssd1 vccd1 vccd1 hold2016/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 _13999_/X vssd1 vssd1 vccd1 vccd1 _17806_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08842_ hold17/X hold83/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08843_/B sky130_fd_sc_hd__mux2_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _17879_/Q vssd1 vssd1 vccd1 vccd1 hold2038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1304 _18226_/Q vssd1 vssd1 vccd1 vccd1 hold1304/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2049 _09103_/X vssd1 vssd1 vccd1 vccd1 _16166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 _18350_/Q vssd1 vssd1 vccd1 vccd1 hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _18220_/Q vssd1 vssd1 vccd1 vccd1 hold1326/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1337 _18209_/Q vssd1 vssd1 vccd1 vccd1 hold1337/X sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ hold8/X hold107/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__mux2_1
Xhold1348 _18298_/Q vssd1 vssd1 vccd1 vccd1 hold1348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _15602_/Q vssd1 vssd1 vccd1 vccd1 hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09325_ _15547_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_164_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ _12813_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _16239_/D sky130_fd_sc_hd__and2_1
XFILLER_0_173_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ _15000_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18042_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09187_ hold1599/X _09218_/B _09186_/X _12789_/A vssd1 vssd1 vccd1 vccd1 _09187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08138_ hold235/X hold369/X hold196/X vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__mux2_1
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ hold2574/X _08082_/B _08068_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08069_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ hold1020/X hold3633/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__mux2_1
X_11080_ hold5441/X _11753_/B _11079_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3240 _16777_/Q vssd1 vssd1 vccd1 vccd1 hold3240/X sky130_fd_sc_hd__dlygate4sd3_1
X_10031_ _16501_/Q _10049_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__and3_1
Xhold3251 _17658_/Q vssd1 vssd1 vccd1 vccd1 hold3251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3262 _10327_/X vssd1 vssd1 vccd1 vccd1 _16599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3273 _17709_/Q vssd1 vssd1 vccd1 vccd1 hold3273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3284 _09649_/X vssd1 vssd1 vccd1 vccd1 _16373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2550 _15722_/Q vssd1 vssd1 vccd1 vccd1 hold2550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3295 _16682_/Q vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2561 _15810_/Q vssd1 vssd1 vccd1 vccd1 hold2561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2572 _15847_/Q vssd1 vssd1 vccd1 vccd1 hold2572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2583 _09097_/X vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2594 _16277_/Q vssd1 vssd1 vccd1 vccd1 hold2594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1860 _08220_/X vssd1 vssd1 vccd1 vccd1 _15746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1871 _14279_/X vssd1 vssd1 vccd1 vccd1 _17940_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14770_ _15217_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14770_/Y sky130_fd_sc_hd__nand2_1
X_11982_ _13749_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__or2_1
Xhold1882 _14091_/X vssd1 vssd1 vccd1 vccd1 _17850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1893 _18316_/Q vssd1 vssd1 vccd1 vccd1 hold1893/X sky130_fd_sc_hd__dlygate4sd3_1
X_13721_ hold2024/X _17694_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ hold4473/X _11222_/B _10932_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _10933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _18353_/CLK _16440_/D vssd1 vssd1 vccd1 vccd1 _16440_/Q sky130_fd_sc_hd__dfxtp_1
X_13652_ hold2820/X _17671_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13653_/B sky130_fd_sc_hd__mux2_1
X_10864_ hold4012/X _11150_/B _10863_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _12909_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _17377_/D sky130_fd_sc_hd__and2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _18386_/CLK _16371_/D vssd1 vssd1 vccd1 vccd1 _16371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13583_ hold2495/X _17648_/Q _13865_/C vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__mux2_1
X_10795_ hold5080/X _11177_/B _10794_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10795_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _18205_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
X_15322_ _15489_/A _15322_/B _15322_/C _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/X
+ sky130_fd_sc_hd__or4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12534_ _12936_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _17354_/D sky130_fd_sc_hd__and2_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _18072_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15253_ _15490_/A1 _15245_/X _15252_/X _15490_/B1 hold3905/X vssd1 vssd1 vccd1 vccd1
+ _15253_/X sky130_fd_sc_hd__a32o_1
X_12465_ hold443/A _12509_/A2 _12505_/A3 _12464_/X _15491_/A vssd1 vssd1 vccd1 vccd1
+ hold347/A sky130_fd_sc_hd__o311a_1
X_14204_ hold730/X _14206_/B vssd1 vssd1 vccd1 vccd1 _14204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11416_ hold4153/X _11792_/B _11415_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15184_ hold1006/X _15219_/B _15183_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15184_/X
+ sky130_fd_sc_hd__o211a_1
X_12396_ _15314_/A _12396_/B vssd1 vssd1 vccd1 vccd1 _17291_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ hold1491/X hold587/X _14134_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14135_/X
+ sky130_fd_sc_hd__o211a_1
X_11347_ hold4611/X _11732_/B _11346_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14066_ _14854_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14066_/X sky130_fd_sc_hd__or2_1
X_11278_ hold5500/X _11762_/B _11277_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _11278_/X
+ sky130_fd_sc_hd__o211a_1
X_10229_ hold2248/X hold3214/X _10523_/S vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__mux2_1
X_13017_ _14980_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__or2_1
X_17825_ _17923_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _18073_/CLK _17756_/D vssd1 vssd1 vccd1 vccd1 _17756_/Q sky130_fd_sc_hd__dfxtp_1
X_14968_ _15129_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__or2_1
X_16707_ _18233_/CLK _16707_/D vssd1 vssd1 vccd1 vccd1 _16707_/Q sky130_fd_sc_hd__dfxtp_1
X_13919_ _14350_/A _13919_/B vssd1 vssd1 vccd1 vccd1 _17767_/D sky130_fd_sc_hd__and2_1
X_17687_ _17719_/CLK _17687_/D vssd1 vssd1 vccd1 vccd1 _17687_/Q sky130_fd_sc_hd__dfxtp_1
X_14899_ hold1932/X hold657/A _14898_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16638_ _18222_/CLK _16638_/D vssd1 vssd1 vccd1 vccd1 _16638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16569_ _18223_/CLK _16569_/D vssd1 vssd1 vccd1 vccd1 _16569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09110_ _15551_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__or2_1
X_18308_ _18308_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09041_ _09047_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _16137_/D sky130_fd_sc_hd__and2_1
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18239_ _18339_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 hold401/A vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 input13/X vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold423 hold423/A vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold434/A vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 hold456/A vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold467 hold467/A vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 data_in[22] vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09943_ hold4885/X _10049_/B _09942_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09943_/X
+ sky130_fd_sc_hd__o211a_1
Xhold489 input63/X vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout903 hold784/X vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__buf_8
Xfanout914 hold770/X vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__buf_8
Xfanout925 hold891/X vssd1 vssd1 vccd1 vccd1 hold756/A sky130_fd_sc_hd__buf_6
Xfanout936 _15207_/A vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__clkbuf_16
X_09874_ hold5189/X _10628_/B _09873_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09874_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout947 _15183_/A vssd1 vssd1 vccd1 vccd1 _15129_/A sky130_fd_sc_hd__buf_8
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _16203_/Q vssd1 vssd1 vccd1 vccd1 hold1101/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _16261_/Q vssd1 vssd1 vccd1 vccd1 hold1112/X sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _09003_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _16031_/D sky130_fd_sc_hd__and2_1
Xhold1123 _13997_/X vssd1 vssd1 vccd1 vccd1 _17805_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _15598_/Q vssd1 vssd1 vccd1 vccd1 hold1134/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 _14243_/X vssd1 vssd1 vccd1 vccd1 _17922_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 hold1339/X vssd1 vssd1 vccd1 vccd1 hold1340/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 _17822_/Q vssd1 vssd1 vccd1 vccd1 hold1167/X sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _15284_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _15998_/D sky130_fd_sc_hd__and2_1
Xhold1178 _08253_/X vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1189 _15787_/Q vssd1 vssd1 vccd1 vccd1 hold1189/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ hold136/X hold426/X _08721_/S vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__mux2_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09308_ hold2370/X _09338_/A2 _09307_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09308_/X
+ sky130_fd_sc_hd__o211a_1
X_10580_ _16684_/Q _10580_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__and3_1
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _15515_/A hold1372/X _09277_/S vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ hold4933/X _13844_/B _12249_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11201_ _16891_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__and3_1
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ hold4536/X _13844_/B _12180_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_249_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17583_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11132_ hold920/X _16868_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _11133_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 hold990/A vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15940_ _17287_/CLK _15940_/D vssd1 vssd1 vccd1 vccd1 hold721/A sky130_fd_sc_hd__dfxtp_1
X_11063_ _18048_/Q hold5608/X _11066_/S vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__mux2_1
Xhold3070 _12695_/X vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10014_ _13150_/A _09918_/A _10013_/X vssd1 vssd1 vccd1 vccd1 _10014_/Y sky130_fd_sc_hd__a21oi_1
Xhold3081 _17390_/Q vssd1 vssd1 vccd1 vccd1 hold3081/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3092 _17405_/Q vssd1 vssd1 vccd1 vccd1 hold3092/X sky130_fd_sc_hd__dlygate4sd3_1
X_15871_ _17742_/CLK _15871_/D vssd1 vssd1 vccd1 vccd1 _15871_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2380 _14769_/X vssd1 vssd1 vccd1 vccd1 _18175_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17610_ _17738_/CLK _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2391 _15130_/X vssd1 vssd1 vccd1 vccd1 _18348_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14822_ _15000_/A _14822_/B vssd1 vssd1 vccd1 vccd1 _14822_/Y sky130_fd_sc_hd__nand2_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _18358_/CLK _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _18323_/Q vssd1 vssd1 vccd1 vccd1 hold1690/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ hold2807/X _14774_/B _14752_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ hold4877/X _12347_/B _11964_/X _08133_/A vssd1 vssd1 vccd1 vccd1 _11965_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _13713_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ _17475_/CLK _17472_/D vssd1 vssd1 vccd1 vccd1 _17472_/Q sky130_fd_sc_hd__dfxtp_1
X_10916_ hold2887/X _16796_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _15185_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__or2_1
X_11896_ hold4389/X _13844_/B _11895_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _11896_/X
+ sky130_fd_sc_hd__o211a_1
X_16423_ _18422_/CLK _16423_/D vssd1 vssd1 vccd1 vccd1 _16423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13734_/A _13635_/B vssd1 vssd1 vccd1 vccd1 _13635_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ hold2853/X _16773_/Q _11153_/C vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16354_ _18395_/CLK _16354_/D vssd1 vssd1 vccd1 vccd1 _16354_/Q sky130_fd_sc_hd__dfxtp_1
X_13566_ _13788_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10778_ hold2501/X _16750_/Q _10874_/S vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ hold632/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12517_ hold1467/X hold3046/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__mux2_1
X_16285_ _18462_/CLK _16285_/D vssd1 vssd1 vccd1 vccd1 _16285_/Q sky130_fd_sc_hd__dfxtp_1
X_13497_ _13791_/A _13497_/B vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18024_ _18035_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
X_15236_ _17327_/Q _09362_/C _15485_/B1 hold84/X vssd1 vssd1 vccd1 vccd1 _15236_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _17317_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _15547_/A hold609/X vssd1 vssd1 vccd1 vccd1 _15167_/Y sky130_fd_sc_hd__nand2_1
X_12379_ _13888_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _14511_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14118_/X sky130_fd_sc_hd__or2_1
X_15098_ hold2816/X _15109_/B _15097_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15098_/X
+ sky130_fd_sc_hd__o211a_1
X_14049_ hold2320/X _14036_/B _14048_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14049_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08610_ _12422_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _15927_/D sky130_fd_sc_hd__and2_1
X_09590_ hold2473/X _13302_/A _10271_/S vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__mux2_1
X_17808_ _17893_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08541_ _15454_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _15894_/D sky130_fd_sc_hd__and2_1
X_17739_ _17739_/CLK _17739_/D vssd1 vssd1 vccd1 vccd1 _17739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08472_ _14866_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08472_/X sky130_fd_sc_hd__or2_1
XFILLER_0_175_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ hold81/X hold727/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5901 _16526_/Q vssd1 vssd1 vccd1 vccd1 hold5901/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5912 _17552_/Q vssd1 vssd1 vccd1 vccd1 hold5912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5923 _17533_/Q vssd1 vssd1 vccd1 vccd1 hold5923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5934 _17556_/Q vssd1 vssd1 vccd1 vccd1 hold5934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5945 hold6005/X vssd1 vssd1 vccd1 vccd1 hold5945/X sky130_fd_sc_hd__buf_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5956 _17943_/Q vssd1 vssd1 vccd1 vccd1 hold5956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5967 _18380_/Q vssd1 vssd1 vccd1 vccd1 hold5967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__clkbuf_4
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5978 _15789_/Q vssd1 vssd1 vccd1 vccd1 hold5978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 input44/X vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5989 data_in[21] vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__buf_8
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _08887_/A vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__clkbuf_4
Xhold297 input58/X vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _08887_/A vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__buf_4
X_09926_ hold3010/X hold5615/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__mux2_1
Xfanout722 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _15032_/A sky130_fd_sc_hd__buf_4
Xfanout733 _15364_/A vssd1 vssd1 vccd1 vccd1 _15052_/A sky130_fd_sc_hd__buf_4
Xfanout744 fanout763/X vssd1 vssd1 vccd1 vccd1 _08111_/A sky130_fd_sc_hd__buf_4
Xfanout755 _14378_/A vssd1 vssd1 vccd1 vccd1 _14380_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout766 _13753_/C1 vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__buf_2
X_09857_ hold1286/X _16443_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__mux2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout777 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _12274_/C1 sky130_fd_sc_hd__buf_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14548_/C1 sky130_fd_sc_hd__buf_4
Xfanout799 fanout816/X vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ hold407/X hold660/X _08864_/S vssd1 vssd1 vccd1 vccd1 hold661/A sky130_fd_sc_hd__mux2_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ hold2816/X hold5681/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__mux2_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ hold32/X hold694/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__mux2_1
XANTENNA_104 _08498_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 hold335/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _15123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _17074_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__and3_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _11097_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__or2_1
XFILLER_0_193_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11681_ hold2170/X hold4538/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__mux2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ hold4836/X _13805_/B _13419_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13420_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10632_ hold3734/X _10542_/A _10631_/X vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13351_ hold4139/X _13829_/B _13350_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10563_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _17258_/Q _12302_/B _13811_/C vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__and3_1
X_16070_ _17307_/CLK _16070_/D vssd1 vssd1 vccd1 vccd1 hold461/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10494_ _10551_/A _10494_/B vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__or2_1
X_13282_ _17586_/Q _17120_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15021_ _15129_/A hold2680/X _15069_/S vssd1 vssd1 vccd1 vccd1 _15022_/B sky130_fd_sc_hd__mux2_1
X_12233_ hold1964/X hold5472/X _12338_/C vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12164_ hold2622/X hold4439/X _12356_/C vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__or2_1
X_12095_ hold2264/X _17189_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__mux2_1
X_16972_ _17852_/CLK _16972_/D vssd1 vssd1 vccd1 vccd1 _16972_/Q sky130_fd_sc_hd__dfxtp_1
X_15923_ _17287_/CLK _15923_/D vssd1 vssd1 vccd1 vccd1 hold697/A sky130_fd_sc_hd__dfxtp_1
X_11046_ _11061_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/X sky130_fd_sc_hd__or2_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _17726_/CLK _15854_/D vssd1 vssd1 vccd1 vccd1 _15854_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ hold1478/X _14822_/B _14804_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14805_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _17748_/CLK _15785_/D vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfxtp_1
X_12997_ hold2945/X _17510_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__mux2_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17524_ _17524_/CLK hold796/X vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _15129_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14736_/X sky130_fd_sc_hd__or2_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11948_ hold1257/X hold3420/X _12332_/C vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17455_ _17456_/CLK _17455_/D vssd1 vssd1 vccd1 vccd1 _17455_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ hold2359/X _14666_/B _14666_/Y _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14667_/X
+ sky130_fd_sc_hd__o211a_1
X_11879_ hold516/X hold3819/X _13871_/C vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__mux2_1
X_16406_ _18319_/CLK _16406_/D vssd1 vssd1 vccd1 vccd1 _16406_/Q sky130_fd_sc_hd__dfxtp_1
X_13618_ hold3498/X _13808_/B _13617_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _13618_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ _18438_/CLK _17386_/D vssd1 vssd1 vccd1 vccd1 _17386_/Q sky130_fd_sc_hd__dfxtp_1
X_14598_ _15099_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ _18378_/CLK _16337_/D vssd1 vssd1 vccd1 vccd1 _16337_/Q sky130_fd_sc_hd__dfxtp_1
X_13549_ hold4850/X _13856_/B _13548_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16268_ _17981_/CLK _16268_/D vssd1 vssd1 vccd1 vccd1 _16268_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5208 _13597_/X vssd1 vssd1 vccd1 vccd1 _17652_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5219 _16012_/Q vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _18071_/CLK hold210/X vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__nand2_1
Xhold4507 _11713_/X vssd1 vssd1 vccd1 vccd1 _17061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4518 _16636_/Q vssd1 vssd1 vccd1 vccd1 hold4518/X sky130_fd_sc_hd__dlygate4sd3_1
X_16199_ _17482_/CLK _16199_/D vssd1 vssd1 vccd1 vccd1 _16199_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4529 _09655_/X vssd1 vssd1 vccd1 vccd1 _16375_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3806 _12321_/Y vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3817 _16487_/Q vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3828 _17121_/Q vssd1 vssd1 vccd1 vccd1 hold3828/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3839 _10062_/Y vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07972_ _15541_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07972_/Y sky130_fd_sc_hd__nand2_1
X_09711_ _11067_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09642_ _09924_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ _10380_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ hold23/X hold599/X _08528_/S vssd1 vssd1 vccd1 vccd1 hold600/A sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ hold2979/X _08488_/B _08454_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08455_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08386_ _14728_/A hold2369/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _09063_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _16120_/D sky130_fd_sc_hd__and2_1
Xhold5720 _10879_/X vssd1 vssd1 vccd1 vccd1 _16783_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5731 _17013_/Q vssd1 vssd1 vccd1 vccd1 hold5731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5742 _10975_/X vssd1 vssd1 vccd1 vccd1 _16815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5753 hold5905/X vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__buf_1
XFILLER_0_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5764 output80/X vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_12
Xhold5775 hold5917/X vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5786 output89/X vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_12
XFILLER_0_130_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5797 hold5927/X vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout530 _09232_/X vssd1 vssd1 vccd1 vccd1 _09277_/S sky130_fd_sc_hd__clkbuf_8
Xfanout541 _12445_/B vssd1 vssd1 vccd1 vccd1 _12505_/A3 sky130_fd_sc_hd__clkbuf_8
X_09909_ _09933_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__or2_1
Xfanout552 _08305_/B vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__clkbuf_8
Xfanout563 _08100_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__clkbuf_8
Xfanout574 _07884_/Y vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__buf_8
Xfanout585 _13244_/S vssd1 vssd1 vccd1 vccd1 _13300_/S sky130_fd_sc_hd__buf_8
X_12920_ hold3269/X _12919_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__mux2_1
Xfanout596 _12910_/S vssd1 vssd1 vccd1 vccd1 _12919_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ hold3225/X _12850_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ hold3871/X _12246_/A _11801_/X vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15570_ _17906_/CLK _15570_/D vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ hold3450/X _12781_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__mux2_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14521_ _14986_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14521_/X sky130_fd_sc_hd__or2_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ hold3759/X _11637_/A _11732_/X vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ _17906_/CLK _17240_/D vssd1 vssd1 vccd1 vccd1 _17240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ hold1399/X _14487_/B _14451_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14452_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11664_ _12246_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ hold2555/X hold4544/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__mux2_1
X_10615_ _10651_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__nor2_1
X_17171_ _17865_/CLK _17171_/D vssd1 vssd1 vccd1 vccd1 _17171_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_264_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17262_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14383_ _14330_/A hold1488/X hold275/X vssd1 vssd1 vccd1 vccd1 _14384_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11595_ _12234_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16122_ _17345_/CLK _16122_/D vssd1 vssd1 vccd1 vccd1 hold388/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ hold2781/X hold3622/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ hold4174/X _10640_/B _10545_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16053_ _17307_/CLK _16053_/D vssd1 vssd1 vccd1 vccd1 _16053_/Q sky130_fd_sc_hd__dfxtp_1
X_13265_ _13265_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__and2_1
X_10477_ hold4105/X _10571_/B _10476_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _10477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15219_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _13794_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13196_ hold5251/X _13195_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_20_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _12255_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__or2_1
X_12078_ _13749_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__or2_1
X_16955_ _17855_/CLK _16955_/D vssd1 vssd1 vccd1 vccd1 _16955_/Q sky130_fd_sc_hd__dfxtp_1
X_15906_ _18425_/CLK _15906_/D vssd1 vssd1 vccd1 vccd1 hold518/A sky130_fd_sc_hd__dfxtp_1
X_11029_ hold4363/X _11222_/B _11028_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _11029_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16886_ _18059_/CLK _16886_/D vssd1 vssd1 vccd1 vccd1 _16886_/Q sky130_fd_sc_hd__dfxtp_1
X_15837_ _17741_/CLK _15837_/D vssd1 vssd1 vccd1 vccd1 _15837_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ _17719_/CLK _15768_/D vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719_ hold2744/X _14718_/B _14718_/Y _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14719_/X
+ sky130_fd_sc_hd__o211a_1
X_17507_ _17517_/CLK _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
X_15699_ _17865_/CLK _15699_/D vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ _14854_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08240_/X sky130_fd_sc_hd__or2_1
X_17438_ _17439_/CLK _17438_/D vssd1 vssd1 vccd1 vccd1 _17438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_26 _15508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_37 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_48 _15515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _15723_/D sky130_fd_sc_hd__and2_1
X_17369_ _17981_/CLK _17369_/D vssd1 vssd1 vccd1 vccd1 _17369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_59 hold29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5005 _16956_/Q vssd1 vssd1 vccd1 vccd1 hold5005/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5016 _12019_/X vssd1 vssd1 vccd1 vccd1 _17163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5027 _11935_/X vssd1 vssd1 vccd1 vccd1 _17135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput100 _13105_/A vssd1 vssd1 vccd1 vccd1 hold5792/A sky130_fd_sc_hd__buf_6
Xhold5038 _16383_/Q vssd1 vssd1 vccd1 vccd1 hold5038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5049 _09871_/X vssd1 vssd1 vccd1 vccd1 _16447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput111 hold5830/X vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_12
Xhold4304 _11632_/X vssd1 vssd1 vccd1 vccd1 _17034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput122 hold5871/X vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_12
Xhold4315 _16650_/Q vssd1 vssd1 vccd1 vccd1 hold4315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4326 _13633_/X vssd1 vssd1 vccd1 vccd1 _17664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput133 hold5846/X vssd1 vssd1 vccd1 vccd1 hold5847/A sky130_fd_sc_hd__buf_6
XFILLER_0_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4337 _16696_/Q vssd1 vssd1 vccd1 vccd1 hold4337/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput144 _13053_/A vssd1 vssd1 vccd1 vccd1 load_status[4] sky130_fd_sc_hd__buf_12
Xhold3603 _11212_/Y vssd1 vssd1 vccd1 vccd1 _16894_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4348 _13738_/X vssd1 vssd1 vccd1 vccd1 _17699_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4359 _16576_/Q vssd1 vssd1 vccd1 vccd1 hold4359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3614 _11784_/Y vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3625 _16530_/Q vssd1 vssd1 vccd1 vccd1 hold3625/X sky130_fd_sc_hd__clkbuf_2
Xhold3636 _16716_/Q vssd1 vssd1 vccd1 vccd1 hold3636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2902 _14761_/X vssd1 vssd1 vccd1 vccd1 _18171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3647 _11749_/Y vssd1 vssd1 vccd1 vccd1 _17073_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2913 _17996_/Q vssd1 vssd1 vccd1 vccd1 hold2913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3658 _15453_/X vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3669 _15423_/X vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 _14921_/X vssd1 vssd1 vccd1 vccd1 _18247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2935 _15514_/X vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07955_ hold1231/X _07991_/A2 _07954_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07955_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2946 _09117_/X vssd1 vssd1 vccd1 vccd1 _16173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2957 _18398_/Q vssd1 vssd1 vccd1 vccd1 hold2957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 _14498_/X vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2979 _15856_/Q vssd1 vssd1 vccd1 vccd1 hold2979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07886_ hold944/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__or2_1
X_09625_ hold3917/X _10001_/B _09624_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _09625_/X
+ sky130_fd_sc_hd__o211a_1
X_09556_ hold4111/X _10571_/B _09555_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _09556_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08507_ hold892/X _08517_/B vssd1 vssd1 vccd1 vccd1 _08507_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09487_ _13056_/C _13030_/A _13034_/D _13053_/A vssd1 vssd1 vccd1 vccd1 _13035_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08438_ hold1328/X _08433_/B _08437_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08369_ _08373_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _15816_/D sky130_fd_sc_hd__and2_1
XFILLER_0_190_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10400_ hold2322/X _16624_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__mux2_1
X_11380_ hold5697/X _11762_/B _11379_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11380_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ hold2793/X hold3342/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5550 _16824_/Q vssd1 vssd1 vccd1 vccd1 hold5550/X sky130_fd_sc_hd__dlygate4sd3_1
X_13050_ _13046_/A _13053_/A _13055_/C vssd1 vssd1 vccd1 vccd1 fanout2/A sky130_fd_sc_hd__a21o_2
X_10262_ hold2955/X hold4224/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10263_/B sky130_fd_sc_hd__mux2_1
Xhold5561 _11296_/X vssd1 vssd1 vccd1 vccd1 _16922_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5572 _16846_/Q vssd1 vssd1 vccd1 vccd1 hold5572/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5583 _10444_/X vssd1 vssd1 vccd1 vccd1 _16638_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12001_ hold4457/X _12308_/B _12000_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5594 _16766_/Q vssd1 vssd1 vccd1 vccd1 hold5594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4860 _17031_/Q vssd1 vssd1 vccd1 vccd1 hold4860/X sky130_fd_sc_hd__dlygate4sd3_1
X_10193_ hold2476/X hold3524/X _10481_/S vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__mux2_1
Xhold4871 _17128_/Q vssd1 vssd1 vccd1 vccd1 hold4871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4882 _11524_/X vssd1 vssd1 vccd1 vccd1 _16998_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4893 _17628_/Q vssd1 vssd1 vccd1 vccd1 hold4893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 _15551_/B vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__clkbuf_4
Xfanout371 _15073_/Y vssd1 vssd1 vccd1 vccd1 _15109_/B sky130_fd_sc_hd__buf_6
Xfanout382 _14842_/Y vssd1 vssd1 vccd1 vccd1 _14880_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16740_ _18071_/CLK _16740_/D vssd1 vssd1 vccd1 vccd1 _16740_/Q sky130_fd_sc_hd__dfxtp_1
X_13952_ _15513_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13952_/X sky130_fd_sc_hd__or2_1
Xfanout393 _14664_/B vssd1 vssd1 vccd1 vccd1 _14666_/B sky130_fd_sc_hd__clkbuf_8
X_12903_ _12909_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _17477_/D sky130_fd_sc_hd__and2_1
X_16671_ _18197_/CLK _16671_/D vssd1 vssd1 vccd1 vccd1 _16671_/Q sky130_fd_sc_hd__dfxtp_1
X_13883_ _17748_/Q _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__and3_1
X_18410_ _18410_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
X_15622_ _17703_/CLK _15622_/D vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _12843_/A _12834_/B vssd1 vssd1 vccd1 vccd1 _17454_/D sky130_fd_sc_hd__and2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18389_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__or2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12765_ _12813_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _17431_/D sky130_fd_sc_hd__and2_1
XFILLER_0_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ hold5960/X _14554_/A2 _14503_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14504_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18272_ _18304_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11716_ hold4852/X _12305_/B _11715_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11716_/X
+ sky130_fd_sc_hd__o211a_1
X_15484_ hold614/X _15484_/A2 _15484_/B1 hold518/X vssd1 vssd1 vccd1 vccd1 _15489_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12849_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _17408_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ _18445_/CLK _17223_/D vssd1 vssd1 vccd1 vccd1 _17223_/Q sky130_fd_sc_hd__dfxtp_1
X_14435_ _15169_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ hold4532/X _12323_/B _11646_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_0_181_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17154_ _17735_/CLK _17154_/D vssd1 vssd1 vccd1 vccd1 _17154_/Q sky130_fd_sc_hd__dfxtp_1
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _15044_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _17982_/D sky130_fd_sc_hd__and2_1
Xinput46 input46/A vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
X_11578_ hold3376/X _11798_/B _11577_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _11578_/X
+ sky130_fd_sc_hd__o211a_1
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
X_16105_ _18405_/CLK _16105_/D vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__dfxtp_1
Xinput68 input68/A vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_13317_ _13800_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _13317_/X sky130_fd_sc_hd__or2_1
Xhold808 hold808/A vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold819 hold819/A vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ hold818/X _16667_/Q _10643_/C vssd1 vssd1 vccd1 vccd1 _10530_/B sky130_fd_sc_hd__mux2_1
X_17085_ _17901_/CLK _17085_/D vssd1 vssd1 vccd1 vccd1 _17085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14297_ hold5964/X _14333_/A2 _14296_/X _14368_/A vssd1 vssd1 vccd1 vccd1 hold625/A
+ sky130_fd_sc_hd__o211a_1
X_16036_ _17292_/CLK _16036_/D vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__dfxtp_1
X_13248_ _13241_/X _13247_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _13178_/X hold5233/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__mux2_1
Xhold2209 next_key vssd1 vssd1 vccd1 vccd1 hold2209/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1508 _09111_/X vssd1 vssd1 vccd1 vccd1 _16170_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ _18052_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 _17987_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1519 _15608_/Q vssd1 vssd1 vccd1 vccd1 hold1519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16938_ _17882_/CLK _16938_/D vssd1 vssd1 vccd1 vccd1 _16938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16869_ _18046_/CLK _16869_/D vssd1 vssd1 vccd1 vccd1 _16869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09410_ _09438_/B _16291_/Q vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _18460_/Q _07802_/B _15490_/A1 vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_133_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_186_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18214_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09272_/A hold144/X vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__and2_1
XFILLER_0_157_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_115_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08223_ _15557_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08154_ _15559_/A hold2195/X hold196/X vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08085_ hold1958/X _08088_/B _08084_/Y _13925_/A vssd1 vssd1 vccd1 vccd1 _08085_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4101 _17041_/Q vssd1 vssd1 vccd1 vccd1 hold4101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4112 _09556_/X vssd1 vssd1 vccd1 vccd1 _16342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4123 _16609_/Q vssd1 vssd1 vccd1 vccd1 hold4123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4134 _11680_/X vssd1 vssd1 vccd1 vccd1 _17050_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3400 _17198_/Q vssd1 vssd1 vccd1 vccd1 hold3400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4145 _16772_/Q vssd1 vssd1 vccd1 vccd1 hold4145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4156 _10294_/X vssd1 vssd1 vccd1 vccd1 _16588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3411 _12701_/X vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3422 _17630_/Q vssd1 vssd1 vccd1 vccd1 hold3422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4167 _17695_/Q vssd1 vssd1 vccd1 vccd1 hold4167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3433 _17032_/Q vssd1 vssd1 vccd1 vccd1 hold3433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4178 _17005_/Q vssd1 vssd1 vccd1 vccd1 hold4178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4189 _10207_/X vssd1 vssd1 vccd1 vccd1 _16559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3444 _17236_/Q vssd1 vssd1 vccd1 vccd1 hold3444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3455 _17435_/Q vssd1 vssd1 vccd1 vccd1 hold3455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2710 _16252_/Q vssd1 vssd1 vccd1 vccd1 hold2710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3466 _17411_/Q vssd1 vssd1 vccd1 vccd1 hold3466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2721 _15663_/Q vssd1 vssd1 vccd1 vccd1 hold2721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2732 _17885_/Q vssd1 vssd1 vccd1 vccd1 hold2732/X sky130_fd_sc_hd__dlygate4sd3_1
X_08987_ hold65/X hold459/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__mux2_1
Xhold3477 _16870_/Q vssd1 vssd1 vccd1 vccd1 hold3477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3488 _10186_/X vssd1 vssd1 vccd1 vccd1 _16552_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _14259_/X vssd1 vssd1 vccd1 vccd1 _17930_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3499 _13618_/X vssd1 vssd1 vccd1 vccd1 _17659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2754 _18060_/Q vssd1 vssd1 vccd1 vccd1 hold2754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2765 _07957_/X vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07938_ _14735_/A _08504_/A vssd1 vssd1 vccd1 vccd1 _07938_/Y sky130_fd_sc_hd__nor2_1
Xhold2776 _18196_/Q vssd1 vssd1 vccd1 vccd1 hold2776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2787 _18255_/Q vssd1 vssd1 vccd1 vccd1 hold2787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2798 _14741_/X vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07869_ _14774_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__nand2_1
X_09608_ hold685/X hold5602/X _11066_/S vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__mux2_1
X_10880_ _17987_/Q _16784_/Q _11171_/C vssd1 vssd1 vccd1 vccd1 _10881_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ hold1432/X _13166_/A _10025_/C vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12550_ hold2447/X _17361_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_148_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ hold2493/X _16991_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ hold184/X _08598_/B _08999_/B _12480_/X _15344_/A vssd1 vssd1 vccd1 vccd1
+ hold185/A sky130_fd_sc_hd__o311a_1
XFILLER_0_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ _14970_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14220_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11432_ hold2607/X _16968_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14151_ hold2038/X _14148_/B _14150_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _14151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ hold1377/X hold4107/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13102_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__or2_1
X_10314_ _10524_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__or2_1
X_14082_ _15535_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14082_/X sky130_fd_sc_hd__or2_1
X_11294_ _17770_/Q hold5289/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5380 _09733_/X vssd1 vssd1 vccd1 vccd1 _16401_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13033_ _13056_/C _13030_/X _13032_/Y vssd1 vssd1 vccd1 vccd1 _13033_/Y sky130_fd_sc_hd__a21oi_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ _18426_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
X_10245_ _10515_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__or2_1
Xhold5391 _16789_/Q vssd1 vssd1 vccd1 vccd1 hold5391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4690 _17040_/Q vssd1 vssd1 vccd1 vccd1 hold4690/X sky130_fd_sc_hd__dlygate4sd3_1
X_10176_ _10380_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
X_17841_ _17873_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14984_ _14984_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__or2_1
X_17772_ _17887_/CLK _17772_/D vssd1 vssd1 vccd1 vccd1 _17772_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout190 fanout209/X vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13935_ _13935_/A hold731/X vssd1 vssd1 vccd1 vccd1 hold732/A sky130_fd_sc_hd__and2_1
X_16723_ _18208_/CLK _16723_/D vssd1 vssd1 vccd1 vccd1 _16723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16654_ _18266_/CLK _16654_/D vssd1 vssd1 vccd1 vccd1 _16654_/Q sky130_fd_sc_hd__dfxtp_1
X_13866_ hold3814/X _13770_/A _13865_/X vssd1 vssd1 vccd1 vccd1 _13866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15605_ _17592_/CLK _15605_/D vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfxtp_1
X_12817_ hold1945/X hold3469/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16585_ _18267_/CLK _16585_/D vssd1 vssd1 vccd1 vccd1 _16585_/Q sky130_fd_sc_hd__dfxtp_1
X_13797_ _13797_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18324_ _18324_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_15536_ hold1760/X _15547_/B _15535_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__o211a_1
X_12748_ _16247_/Q hold3025/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux2_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18255_ _18319_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ hold493/X _09365_/B _09362_/D hold327/X vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__a22o_1
X_12679_ _18455_/Q _17404_/Q _12679_/S vssd1 vssd1 vccd1 vccd1 _12679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _17906_/CLK _17206_/D vssd1 vssd1 vccd1 vccd1 _17206_/Q sky130_fd_sc_hd__dfxtp_1
X_14418_ hold5963/X hold209/X _14417_/X _14418_/C1 vssd1 vssd1 vccd1 vccd1 hold210/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18186_ _18218_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ hold421/X _09386_/A _09392_/D hold395/X vssd1 vssd1 vccd1 vccd1 _15398_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17137_ _17900_/CLK _17137_/D vssd1 vssd1 vccd1 vccd1 _17137_/Q sky130_fd_sc_hd__dfxtp_1
X_14349_ _15191_/A hold1171/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__mux2_1
Xhold605 input57/X vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__buf_1
XFILLER_0_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold616 hold628/X vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__clkbuf_4
Xhold627 hold627/A vssd1 vssd1 vccd1 vccd1 input70/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 hold649/A vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ _17852_/CLK _17068_/D vssd1 vssd1 vccd1 vccd1 _17068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _17528_/CLK _16019_/D vssd1 vssd1 vccd1 vccd1 hold707/A sky130_fd_sc_hd__dfxtp_1
X_08910_ hold5/X hold259/X _08910_/S vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ hold1962/X _16454_/Q _11201_/C vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__mux2_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _15870_/Q vssd1 vssd1 vccd1 vccd1 hold2006/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2017 _14889_/X vssd1 vssd1 vccd1 vccd1 _18233_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08841_ _15394_/A _08841_/B vssd1 vssd1 vccd1 vccd1 _16039_/D sky130_fd_sc_hd__and2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _15792_/Q vssd1 vssd1 vccd1 vccd1 hold2028/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 _14151_/X vssd1 vssd1 vccd1 vccd1 _17879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1305 _14875_/X vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _15134_/X vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1327 _14863_/X vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ _08970_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _16006_/D sky130_fd_sc_hd__and2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 _14839_/X vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1349 _17831_/Q vssd1 vssd1 vccd1 vccd1 hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ hold2165/X _09325_/B _09323_/Y _15506_/A vssd1 vssd1 vccd1 vccd1 _09324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _15531_/A hold1081/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08206_ hold1218/X _08209_/B _08205_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08206_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ _15515_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08137_ _08137_/A _08137_/B vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08068_ _15527_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18438_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3230 _17159_/Q vssd1 vssd1 vccd1 vccd1 hold3230/X sky130_fd_sc_hd__dlygate4sd3_1
X_10030_ _10588_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__nor2_1
Xhold3241 _10765_/X vssd1 vssd1 vccd1 vccd1 _16745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3252 _13519_/X vssd1 vssd1 vccd1 vccd1 _17626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3263 _16436_/Q vssd1 vssd1 vccd1 vccd1 hold3263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3274 _13672_/X vssd1 vssd1 vccd1 vccd1 _17677_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2540 _16228_/Q vssd1 vssd1 vccd1 vccd1 hold2540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3285 _16472_/Q vssd1 vssd1 vccd1 vccd1 hold3285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2551 _17865_/Q vssd1 vssd1 vccd1 vccd1 hold2551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3296 _10480_/X vssd1 vssd1 vccd1 vccd1 _16650_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2562 _15836_/Q vssd1 vssd1 vccd1 vccd1 hold2562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2573 _08434_/X vssd1 vssd1 vccd1 vccd1 _15847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2584 _18207_/Q vssd1 vssd1 vccd1 vccd1 hold2584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1850 _15768_/Q vssd1 vssd1 vccd1 vccd1 hold1850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 _09334_/X vssd1 vssd1 vccd1 vccd1 _16277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1861 _15632_/Q vssd1 vssd1 vccd1 vccd1 hold1861/X sky130_fd_sc_hd__dlygate4sd3_1
X_11981_ hold1395/X hold3370/X _13844_/C vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__mux2_1
Xhold1872 _17917_/Q vssd1 vssd1 vccd1 vccd1 hold1872/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1883 _17516_/Q vssd1 vssd1 vccd1 vccd1 hold1883/X sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ hold4331/X _13814_/B _13719_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13720_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1894 _16271_/Q vssd1 vssd1 vccd1 vccd1 hold1894/X sky130_fd_sc_hd__dlygate4sd3_1
X_10932_ _11031_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10932_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ hold4844/X _13859_/B _13650_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13651_/X
+ sky130_fd_sc_hd__o211a_1
X_10863_ _11061_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ hold3008/X _12601_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16370_ _18315_/CLK _16370_/D vssd1 vssd1 vccd1 vccd1 _16370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13582_ hold3556/X _13847_/B _13581_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13582_/X
+ sky130_fd_sc_hd__o211a_1
X_10794_ _11082_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__or2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15321_ _16296_/Q _15477_/A2 _15487_/B1 hold394/X _15320_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ hold3438/X _12532_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__mux2_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _18046_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
X_15252_ _15489_/A _15252_/B _15252_/C _15252_/D vssd1 vssd1 vccd1 vccd1 _15252_/X
+ sky130_fd_sc_hd__or4_1
X_12464_ _17325_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ hold2270/X _14202_/B _14202_/Y _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14203_/X
+ sky130_fd_sc_hd__o211a_1
X_11415_ _11697_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__or2_1
X_15183_ _15183_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12395_ hold47/X hold560/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ _15207_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14134_/X sky130_fd_sc_hd__or2_1
X_11346_ _11637_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ hold991/X _14105_/A2 _14064_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 hold992/A
+ sky130_fd_sc_hd__o211a_1
X_11277_ _11667_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11277_/X sky130_fd_sc_hd__or2_1
X_13016_ hold1883/X _13003_/Y _13015_/X _12936_/A vssd1 vssd1 vccd1 vccd1 _13016_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10228_ hold4459/X _10646_/B _10227_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _17855_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_1
X_10159_ hold4453/X _10619_/B _10158_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10159_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17755_ _18009_/CLK _17755_/D vssd1 vssd1 vccd1 vccd1 _17755_/Q sky130_fd_sc_hd__dfxtp_1
X_14967_ _15508_/A hold656/X vssd1 vssd1 vccd1 vccd1 _15012_/B sky130_fd_sc_hd__or2_4
X_16706_ _18220_/CLK _16706_/D vssd1 vssd1 vccd1 vccd1 _16706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ _15207_/A hold1319/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__mux2_1
X_17686_ _17686_/CLK _17686_/D vssd1 vssd1 vccd1 vccd1 _17686_/Q sky130_fd_sc_hd__dfxtp_1
X_14898_ _15129_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16637_ _18219_/CLK _16637_/D vssd1 vssd1 vccd1 vccd1 _16637_/Q sky130_fd_sc_hd__dfxtp_1
X_13849_ _13873_/A _13849_/B vssd1 vssd1 vccd1 vccd1 _13849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16568_ _18126_/CLK _16568_/D vssd1 vssd1 vccd1 vccd1 _16568_/Q sky130_fd_sc_hd__dfxtp_1
X_18307_ _18371_/CLK hold131/X vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
X_15519_ _15519_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__or2_1
X_16499_ _18386_/CLK _16499_/D vssd1 vssd1 vccd1 vccd1 _16499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09040_ hold5/X hold112/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ _18398_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18169_ _18230_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold402 hold402/A vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold413/A vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 hold446/A vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 hold468/A vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _09954_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__or2_1
Xhold479 hold479/A vssd1 vssd1 vccd1 vccd1 input19/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout904 hold784/X vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__clkbuf_4
Xfanout915 hold770/X vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__clkbuf_4
Xfanout926 hold891/X vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__buf_4
X_09873_ _10491_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__or2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 _15207_/A vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__clkbuf_16
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 hold943/X vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__clkbuf_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ hold53/X hold538/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__mux2_1
Xhold1102 _09183_/X vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _09302_/X vssd1 vssd1 vccd1 vccd1 _16261_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _18045_/Q vssd1 vssd1 vccd1 vccd1 hold1124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _07909_/X vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 _15878_/Q vssd1 vssd1 vccd1 vccd1 hold1146/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ hold81/X hold506/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08756_/B sky130_fd_sc_hd__mux2_1
Xhold1157 hold1341/X vssd1 vssd1 vccd1 vccd1 hold1157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _14033_/X vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _16206_/Q vssd1 vssd1 vccd1 vccd1 hold1179/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _15491_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _15964_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_130_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09307_ _14988_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ _12789_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _16230_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09169_ hold1381/X _09164_/B _09168_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _11218_/A _11200_/B vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12180_ _13749_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ hold5672/X _11765_/B _11130_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11131_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ hold4043/X _11150_/B _11061_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _11062_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_289_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3060 _18301_/Q vssd1 vssd1 vccd1 vccd1 hold3060/X sky130_fd_sc_hd__dlygate4sd3_1
X_10013_ _16495_/Q _10013_/B _10028_/C vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__and3_1
Xhold3071 _17370_/Q vssd1 vssd1 vccd1 vccd1 hold3071/X sky130_fd_sc_hd__dlygate4sd3_1
X_15870_ _17678_/CLK _15870_/D vssd1 vssd1 vccd1 vccd1 _15870_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3082 _12641_/X vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3093 _17393_/Q vssd1 vssd1 vccd1 vccd1 hold3093/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_218_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17895_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2370 _16264_/Q vssd1 vssd1 vccd1 vccd1 hold2370/X sky130_fd_sc_hd__dlygate4sd3_1
X_14821_ hold1110/X _14822_/B _14820_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14821_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2381 _18347_/Q vssd1 vssd1 vccd1 vccd1 hold2381/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2392 _15635_/Q vssd1 vssd1 vccd1 vccd1 hold2392/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1680 _13955_/X vssd1 vssd1 vccd1 vccd1 _17784_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17540_ _18386_/CLK _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1691 _15078_/X vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14752_ _14984_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12255_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__or2_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ hold1807/X _17688_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__mux2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _18451_/CLK _17471_/D vssd1 vssd1 vccd1 vccd1 _17471_/Q sky130_fd_sc_hd__dfxtp_1
X_10915_ hold4186/X _11201_/B _10914_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _10915_/X
+ sky130_fd_sc_hd__o211a_1
X_14683_ hold2685/X _14718_/B _14682_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14683_/X
+ sky130_fd_sc_hd__o211a_1
X_11895_ _13749_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__or2_1
X_13634_ hold2199/X _17665_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__mux2_1
X_16422_ _18337_/CLK _16422_/D vssd1 vssd1 vccd1 vccd1 _16422_/Q sky130_fd_sc_hd__dfxtp_1
X_10846_ hold4257/X _11735_/B _10845_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _10846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ _18330_/CLK _16353_/D vssd1 vssd1 vccd1 vccd1 _16353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13565_ hold2108/X hold5179/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13566_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ hold4587/X _11735_/B _10776_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _10777_/X
+ sky130_fd_sc_hd__o211a_1
X_15304_ _15304_/A _15304_/B vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12516_ _13002_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _17348_/D sky130_fd_sc_hd__and2_1
X_16284_ _18243_/CLK _16284_/D vssd1 vssd1 vccd1 vccd1 _16284_/Q sky130_fd_sc_hd__dfxtp_1
X_13496_ hold2679/X hold5060/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13497_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15235_ _15993_/Q _15483_/B vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__or2_1
X_18023_ _18055_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ hold23/X _08598_/B _08999_/B _12446_/X _09047_/A vssd1 vssd1 vccd1 vccd1
+ hold24/A sky130_fd_sc_hd__o311a_1
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ hold2478/X hold609/X _15165_/Y _15060_/A vssd1 vssd1 vccd1 vccd1 _15166_/X
+ sky130_fd_sc_hd__o211a_1
X_12378_ hold3767/X _12282_/A _12377_/X vssd1 vssd1 vccd1 vccd1 _12378_/Y sky130_fd_sc_hd__a21oi_1
X_14117_ hold1544/X hold587/X _14116_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _14117_/X
+ sky130_fd_sc_hd__o211a_1
X_11329_ hold4854/X _12305_/B _11328_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15097_ _15205_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _14728_/A _14050_/B vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17807_ _17829_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_1
X_15999_ _18406_/CLK _15999_/D vssd1 vssd1 vccd1 vccd1 hold706/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08540_ hold32/X hold703/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17738_ _17738_/CLK _17738_/D vssd1 vssd1 vccd1 vccd1 _17738_/Q sky130_fd_sc_hd__dfxtp_1
X_08471_ hold908/X _08486_/B _08470_/X _08151_/A vssd1 vssd1 vccd1 vccd1 hold909/A
+ sky130_fd_sc_hd__o211a_1
X_17669_ _17669_/CLK _17669_/D vssd1 vssd1 vccd1 vccd1 _17669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09023_ _09063_/A hold526/X vssd1 vssd1 vccd1 vccd1 _16128_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5902 _16929_/Q vssd1 vssd1 vccd1 vccd1 hold5902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5913 _17547_/Q vssd1 vssd1 vccd1 vccd1 hold5913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5924 _17553_/Q vssd1 vssd1 vccd1 vccd1 hold5924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5935 _17526_/Q vssd1 vssd1 vccd1 vccd1 hold5935/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5946 data_in[2] vssd1 vssd1 vccd1 vccd1 hold404/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 la_data_in[17] vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5957 _18187_/Q vssd1 vssd1 vccd1 vccd1 hold5957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__buf_1
Xhold5968 _17914_/Q vssd1 vssd1 vccd1 vccd1 hold5968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold40/X vssd1 vssd1 vccd1 vccd1 input32/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5979 _18018_/Q vssd1 vssd1 vccd1 vccd1 hold5979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__buf_4
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _08887_/A vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__clkbuf_2
X_09925_ hold5383/X _10025_/B _09924_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09925_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout712 _08585_/A vssd1 vssd1 vccd1 vccd1 _08887_/A sky130_fd_sc_hd__clkbuf_4
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout723 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _15038_/A sky130_fd_sc_hd__buf_2
Xfanout734 _14985_/C1 vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__buf_2
Xfanout745 _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__buf_4
Xfanout756 fanout763/X vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__buf_2
X_09856_ hold5072/X _09952_/A2 _09855_/X _15144_/C1 vssd1 vssd1 vccd1 vccd1 _09856_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout767 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _13753_/C1 sky130_fd_sc_hd__buf_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_311_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17128_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout778 _14191_/C1 vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__buf_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 _08257_/C1 vssd1 vssd1 vccd1 vccd1 _14546_/C1 sky130_fd_sc_hd__clkbuf_4
X_08807_ _09003_/A _08807_/B vssd1 vssd1 vccd1 vccd1 _16022_/D sky130_fd_sc_hd__and2_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ hold5098/X _10073_/B _09786_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09787_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _09003_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _15989_/D sky130_fd_sc_hd__and2_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 fanout337/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 hold335/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ hold407/X hold416/X _08669_/S vssd1 vssd1 vccd1 vccd1 hold417/A sky130_fd_sc_hd__mux2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ hold2899/X hold3849/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11680_ _11774_/A _11783_/B _11679_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11680_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _16701_/Q _10631_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10631_/X sky130_fd_sc_hd__and3_1
XFILLER_0_107_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _13734_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ hold2703/X hold3531/X _10562_/S vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ _12301_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _12301_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _13281_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__and2_1
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ hold1324/X hold4157/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ hold300/X hold656/A vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__or2_1
X_12232_ hold4903/X _12362_/B _12231_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12163_ hold4981/X _12311_/B _12162_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _12163_/X
+ sky130_fd_sc_hd__o211a_1
X_11114_ hold2012/X _16862_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12094_ hold4729/X _12320_/B _12093_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _12094_/X
+ sky130_fd_sc_hd__o211a_1
X_16971_ _17884_/CLK _16971_/D vssd1 vssd1 vccd1 vccd1 _16971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15922_ _18408_/CLK _15922_/D vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__dfxtp_1
X_11045_ hold2246/X _16839_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _17742_/CLK _15853_/D vssd1 vssd1 vccd1 vccd1 _15853_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _15197_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__or2_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15784_ _17737_/CLK _15784_/D vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfxtp_1
X_12996_ _12996_/A _12996_/B vssd1 vssd1 vccd1 vccd1 _17508_/D sky130_fd_sc_hd__and2_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _17523_/CLK _17523_/D vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ hold5375/X _12329_/B _11946_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11947_/X
+ sky130_fd_sc_hd__o211a_1
X_14735_ _14735_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14784_/B sky130_fd_sc_hd__or2_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _18456_/CLK _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14666_ _14774_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14666_/Y sky130_fd_sc_hd__nand2_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ hold4597/X _12356_/B _11877_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _11878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16405_ _18382_/CLK _16405_/D vssd1 vssd1 vccd1 vccd1 _16405_/Q sky130_fd_sc_hd__dfxtp_1
X_13617_ _13713_/A _13617_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__or2_1
X_10829_ hold2489/X _16767_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__mux2_1
X_17385_ _18438_/CLK _17385_/D vssd1 vssd1 vccd1 vccd1 _17385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ hold2884/X _14612_/B _14596_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13548_ _13776_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__or2_1
X_16336_ _18385_/CLK _16336_/D vssd1 vssd1 vccd1 vccd1 _16336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16267_ _17496_/CLK _16267_/D vssd1 vssd1 vccd1 vccd1 _16267_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ _13737_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__or2_1
Xhold5209 _17748_/Q vssd1 vssd1 vccd1 vccd1 hold5209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _18069_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
X_15218_ hold2002/X _15221_/B _15217_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 _15218_/X
+ sky130_fd_sc_hd__o211a_1
X_16198_ _17475_/CLK _16198_/D vssd1 vssd1 vccd1 vccd1 _16198_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4508 _16987_/Q vssd1 vssd1 vccd1 vccd1 hold4508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4519 _10342_/X vssd1 vssd1 vccd1 vccd1 _16604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ hold747/X _15149_/B vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__or2_1
Xhold3807 _12322_/Y vssd1 vssd1 vccd1 vccd1 _17264_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3818 _09895_/X vssd1 vssd1 vccd1 vccd1 _16455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3829 _12372_/Y vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07971_ hold1375/X _07978_/B _07970_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _07971_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ _18307_/Q _16394_/Q _11066_/S vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__mux2_1
X_09641_ hold2234/X _16371_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09572_ hold865/X _13254_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ _08730_/A _13046_/C vssd1 vssd1 vccd1 vccd1 _08528_/S sky130_fd_sc_hd__or2_2
XFILLER_0_136_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08454_ _15513_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08454_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _08389_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _15824_/D sky130_fd_sc_hd__and2_1
XFILLER_0_175_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ hold35/X hold476/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5710 _11407_/X vssd1 vssd1 vccd1 vccd1 _16959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5721 _17047_/Q vssd1 vssd1 vccd1 vccd1 hold5721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5732 _11473_/X vssd1 vssd1 vccd1 vccd1 _16981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5743 _17055_/Q vssd1 vssd1 vccd1 vccd1 hold5743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5754 output83/X vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5765 hold5911/X vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__buf_1
Xhold5776 output77/X vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_12
Xhold5787 hold5921/X vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5798 output92/X vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_12
XFILLER_0_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout520 _10523_/S vssd1 vssd1 vccd1 vccd1 _10619_/C sky130_fd_sc_hd__clkbuf_8
Xfanout531 _09228_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__buf_4
Xfanout542 _08860_/S vssd1 vssd1 vccd1 vccd1 _08864_/S sky130_fd_sc_hd__buf_8
X_09908_ hold2459/X hold5399/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__mux2_1
Xfanout553 _08336_/A2 vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__clkbuf_8
Xfanout564 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__buf_8
Xfanout575 _07873_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__clkbuf_8
Xfanout586 _13308_/S vssd1 vssd1 vccd1 vccd1 _13244_/S sky130_fd_sc_hd__buf_8
X_09839_ hold1315/X hold5350/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout597 _12910_/S vssd1 vssd1 vccd1 vccd1 _12922_/S sky130_fd_sc_hd__clkbuf_8
X_12850_ hold973/X hold3199/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _17091_/Q _12341_/B _12341_/C vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__and3_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ hold1179/X hold3048/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__mux2_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ hold2862/X _14554_/A2 _14519_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14520_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _17068_/Q _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__and3_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14451_ hold756/X _14499_/B vssd1 vssd1 vccd1 vccd1 _14451_/X sky130_fd_sc_hd__or2_1
X_11663_ hold1204/X hold4121/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ hold5060/X _13880_/B _13401_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13402_/X
+ sky130_fd_sc_hd__o211a_1
X_10614_ hold3628/X _10422_/A _10613_/X vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17170_ _17170_/CLK _17170_/D vssd1 vssd1 vccd1 vccd1 _17170_/Q sky130_fd_sc_hd__dfxtp_1
X_14382_ _14382_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__and2_1
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ hold1249/X _17022_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__mux2_1
X_16121_ _17522_/CLK _16121_/D vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ hold4828/X _13811_/B _13332_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10545_ _10554_/A _10545_/B vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _17343_/CLK _16052_/D vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__dfxtp_1
X_13264_ _13257_/X _13263_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ _10560_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15003_ hold867/X _15006_/B _15002_/Y _15003_/C1 vssd1 vssd1 vccd1 vccd1 hold868/A
+ sky130_fd_sc_hd__o211a_1
X_12215_ hold2334/X _17229_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12216_/B sky130_fd_sc_hd__mux2_1
X_13195_ _13194_/X _16917_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_233_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17216_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12146_ hold1694/X _17206_/Q _13388_/S vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ hold2836/X hold4335/X _13844_/C vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__mux2_1
X_16954_ _17894_/CLK _16954_/D vssd1 vssd1 vccd1 vccd1 _16954_/Q sky130_fd_sc_hd__dfxtp_1
X_15905_ _17300_/CLK _15905_/D vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__dfxtp_1
X_11028_ _11031_/A _11028_/B vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__or2_1
X_16885_ _18066_/CLK _16885_/D vssd1 vssd1 vccd1 vccd1 _16885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _17697_/CLK _15836_/D vssd1 vssd1 vccd1 vccd1 _15836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _17686_/CLK _15767_/D vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfxtp_1
X_12979_ hold2374/X _17504_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__mux2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ _17506_/CLK _17506_/D vssd1 vssd1 vccd1 vccd1 _17506_/Q sky130_fd_sc_hd__dfxtp_1
X_14718_ _15219_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15698_ _17268_/CLK _15698_/D vssd1 vssd1 vccd1 vccd1 _15698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17437_ _17439_/CLK _17437_/D vssd1 vssd1 vccd1 vccd1 _17437_/Q sky130_fd_sc_hd__dfxtp_1
X_14649_ hold2187/X _14664_/B _14648_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14649_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_27 _15508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _15521_/A hold2813/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17368_ _17496_/CLK _17368_/D vssd1 vssd1 vccd1 vccd1 _17368_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_49 _15515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _18460_/CLK _16319_/D vssd1 vssd1 vccd1 vccd1 _16319_/Q sky130_fd_sc_hd__dfxtp_1
X_17299_ _18411_/CLK _17299_/D vssd1 vssd1 vccd1 vccd1 hold596/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5006 _11302_/X vssd1 vssd1 vccd1 vccd1 _16924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5017 _16410_/Q vssd1 vssd1 vccd1 vccd1 hold5017/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5028 _17131_/Q vssd1 vssd1 vccd1 vccd1 hold5028/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput101 _13113_/A vssd1 vssd1 vccd1 vccd1 hold5790/A sky130_fd_sc_hd__buf_6
Xhold5039 _09583_/X vssd1 vssd1 vccd1 vccd1 _16351_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4305 _16607_/Q vssd1 vssd1 vccd1 vccd1 hold4305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 hold5181/X vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_12
Xoutput123 hold5862/X vssd1 vssd1 vccd1 vccd1 hold5863/A sky130_fd_sc_hd__buf_6
Xhold4316 _10384_/X vssd1 vssd1 vccd1 vccd1 _16618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4327 _16637_/Q vssd1 vssd1 vccd1 vccd1 hold4327/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput134 hold5841/X vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_12
Xoutput145 _13046_/A vssd1 vssd1 vccd1 vccd1 load_status[5] sky130_fd_sc_hd__buf_12
Xhold4338 _10522_/X vssd1 vssd1 vccd1 vccd1 _16664_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4349 _16559_/Q vssd1 vssd1 vccd1 vccd1 hold4349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3604 _16719_/Q vssd1 vssd1 vccd1 vccd1 hold3604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3615 _11785_/Y vssd1 vssd1 vccd1 vccd1 _17085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3626 _10599_/Y vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3637 _11157_/Y vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2903 _18025_/Q vssd1 vssd1 vccd1 vccd1 hold2903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3648 _16723_/Q vssd1 vssd1 vccd1 vccd1 hold3648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3659 _16348_/Q vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2914 _14396_/X vssd1 vssd1 vccd1 vccd1 _17996_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2925 _17371_/Q vssd1 vssd1 vccd1 vccd1 hold2925/X sky130_fd_sc_hd__dlygate4sd3_1
X_07954_ _14517_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2936 _17921_/Q vssd1 vssd1 vccd1 vccd1 hold2936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2947 _18001_/Q vssd1 vssd1 vccd1 vccd1 hold2947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2958 _15232_/X vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2969 _18072_/Q vssd1 vssd1 vccd1 vccd1 hold2969/X sky130_fd_sc_hd__dlygate4sd3_1
X_07885_ hold816/X hold585/X vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__or2_4
X_09624_ _09948_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09555_ _10380_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17984_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08506_ hold1788/X _08503_/Y _08505_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _08506_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09486_ hold1601/X hold5887/X _09485_/Y vssd1 vssd1 vccd1 vccd1 _16323_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08437_ _14330_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08368_ _15537_/A hold1929/X hold122/X vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08299_ _14517_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08299_/X sky130_fd_sc_hd__or2_1
X_10330_ hold3936/X _10897_/A2 _10329_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _10330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5540 _17018_/Q vssd1 vssd1 vccd1 vccd1 hold5540/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5551 _10906_/X vssd1 vssd1 vccd1 vccd1 _16792_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10261_ hold4123/X _10643_/B _10260_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5562 _16391_/Q vssd1 vssd1 vccd1 vccd1 hold5562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5573 _10972_/X vssd1 vssd1 vccd1 vccd1 _16814_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12000_ _13797_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__or2_1
Xhold5584 _16856_/Q vssd1 vssd1 vccd1 vccd1 hold5584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4850 _17668_/Q vssd1 vssd1 vccd1 vccd1 hold4850/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5595 _10732_/X vssd1 vssd1 vccd1 vccd1 _16734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4861 _11527_/X vssd1 vssd1 vccd1 vccd1 _16999_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10192_ hold3533/X _10558_/A2 _10191_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _10192_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4872 _11818_/X vssd1 vssd1 vccd1 vccd1 _17096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4883 _16615_/Q vssd1 vssd1 vccd1 vccd1 hold4883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4894 _13429_/X vssd1 vssd1 vccd1 vccd1 _17596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout350 _08930_/S vssd1 vssd1 vccd1 vccd1 _08932_/S sky130_fd_sc_hd__buf_6
Xfanout361 _15560_/A2 vssd1 vssd1 vccd1 vccd1 _15547_/B sky130_fd_sc_hd__buf_4
XFILLER_0_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout372 hold301/X vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__buf_6
X_13951_ hold1229/X _13980_/B _13950_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _13951_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout383 _14838_/B vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__buf_6
Xfanout394 _14626_/Y vssd1 vssd1 vccd1 vccd1 _14664_/B sky130_fd_sc_hd__buf_6
X_12902_ hold3004/X _12901_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__mux2_1
X_13882_ _13888_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13882_/Y sky130_fd_sc_hd__nor2_1
X_16670_ _18228_/CLK _16670_/D vssd1 vssd1 vccd1 vccd1 _16670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15621_ _17217_/CLK _15621_/D vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfxtp_1
X_12833_ hold3091/X _12832_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__mux2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18340_ _18380_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ hold3541/X _12763_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__mux2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ hold1223/X _15547_/B _15551_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _15552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _12018_/A _11715_/B vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__or2_1
X_14503_ _15183_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__or2_1
X_15483_ hold599/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__or2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _18337_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
X_12695_ hold3069/X _12694_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__mux2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17222_ _17719_/CLK _17222_/D vssd1 vssd1 vccd1 vccd1 _17222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11646_ _12036_/A _11646_/B vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__or2_1
X_14434_ hold2094/X _14433_/B _14433_/Y _14368_/A vssd1 vssd1 vccd1 vccd1 _14434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 input14/A vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput25 input25/A vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17153_ _17217_/CLK _17153_/D vssd1 vssd1 vccd1 vccd1 _17153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14365_ _15099_/A hold2490/X hold275/X vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__mux2_1
Xinput36 input36/A vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ _11697_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__or2_1
Xinput47 input47/A vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
X_16104_ _18417_/CLK _16104_/D vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dfxtp_1
X_13316_ hold962/X _17559_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__mux2_1
Xinput58 input58/A vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
Xinput69 input69/A vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
X_10528_ hold4575/X _10640_/B _10527_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10528_/X
+ sky130_fd_sc_hd__o211a_1
X_17084_ _17900_/CLK _17084_/D vssd1 vssd1 vccd1 vccd1 _17084_/Q sky130_fd_sc_hd__dfxtp_1
Xhold809 hold809/A vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ hold490/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _13311_/A1 _13245_/X _13246_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13247_/X
+ sky130_fd_sc_hd__o211a_1
X_16035_ _18407_/CLK _16035_/D vssd1 vssd1 vccd1 vccd1 hold648/A sky130_fd_sc_hd__dfxtp_1
X_10459_ hold3221/X _10649_/B _10458_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10459_/X
+ sky130_fd_sc_hd__o211a_1
X_13178_ _17573_/Q _17107_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__mux2_1
X_12129_ _13794_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or2_1
X_17986_ _18062_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__dfxtp_1
Xhold1509 _15771_/Q vssd1 vssd1 vccd1 vccd1 hold1509/X sky130_fd_sc_hd__dlygate4sd3_1
X_16937_ _17785_/CLK _16937_/D vssd1 vssd1 vccd1 vccd1 _16937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16868_ _18071_/CLK _16868_/D vssd1 vssd1 vccd1 vccd1 _16868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15819_ _17634_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 _15819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16799_ _18034_/CLK _16799_/D vssd1 vssd1 vccd1 vccd1 _16799_/Q sky130_fd_sc_hd__dfxtp_1
X_09340_ _18460_/Q _07802_/B _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ hold173/A _16247_/Q _09277_/S vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ hold2639/X _08209_/B _08221_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _08222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_155_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18219_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08084_ _15217_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_141_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4102 _11557_/X vssd1 vssd1 vccd1 vccd1 _17009_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4113 _17050_/Q vssd1 vssd1 vccd1 vccd1 hold4113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4124 _10261_/X vssd1 vssd1 vccd1 vccd1 _16577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4135 _17624_/Q vssd1 vssd1 vccd1 vccd1 hold4135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3401 _12028_/X vssd1 vssd1 vccd1 vccd1 _17166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4146 _10750_/X vssd1 vssd1 vccd1 vccd1 _16740_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4157 _16655_/Q vssd1 vssd1 vccd1 vccd1 hold4157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3412 _17409_/Q vssd1 vssd1 vccd1 vccd1 hold3412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3423 _13435_/X vssd1 vssd1 vccd1 vccd1 _17598_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4168 _13630_/X vssd1 vssd1 vccd1 vccd1 _17663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3434 _11530_/X vssd1 vssd1 vccd1 vccd1 _17000_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4179 _11449_/X vssd1 vssd1 vccd1 vccd1 _16973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3445 _12142_/X vssd1 vssd1 vccd1 vccd1 _17204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2700 _14239_/X vssd1 vssd1 vccd1 vccd1 _17920_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2711 _18281_/Q vssd1 vssd1 vccd1 vccd1 hold2711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3456 _17509_/Q vssd1 vssd1 vccd1 vccd1 hold3456/X sky130_fd_sc_hd__dlygate4sd3_1
X_08986_ _15344_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _16110_/D sky130_fd_sc_hd__and2_1
Xhold2722 _08044_/X vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3467 _17510_/Q vssd1 vssd1 vccd1 vccd1 hold3467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2733 _14165_/X vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3478 _11044_/X vssd1 vssd1 vccd1 vccd1 _16838_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2744 _18151_/Q vssd1 vssd1 vccd1 vccd1 hold2744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3489 _17416_/Q vssd1 vssd1 vccd1 vccd1 hold3489/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2755 _14528_/X vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07937_ hold2388/X _07924_/B _07936_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _07937_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2766 _15697_/Q vssd1 vssd1 vccd1 vccd1 hold2766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2777 _14813_/X vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2788 _14937_/X vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 _18183_/Q vssd1 vssd1 vccd1 vccd1 hold2799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07868_ hold2129/X _07869_/B _07867_/Y _12256_/C1 vssd1 vssd1 vccd1 vccd1 _07868_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09607_ hold5562/X _09998_/B _09606_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07799_ _11155_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ hold5699/X _10016_/B _09537_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09472_/B _09472_/C _09472_/D vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__and3_1
X_11500_ hold5466/X _12329_/B _11499_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11500_/X
+ sky130_fd_sc_hd__o211a_1
X_12480_ _17333_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ hold4700/X _12299_/B _11430_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11431_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14150_ _15549_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14150_/X sky130_fd_sc_hd__or2_1
X_11362_ hold4441/X _12320_/B _11361_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11362_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13101_ _13100_/X hold3662/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__mux2_1
X_10313_ hold1952/X _16595_/Q _10619_/C vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ hold2509/X _14094_/B _14080_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14081_/X
+ sky130_fd_sc_hd__o211a_1
X_11293_ hold5443/X _12338_/B _11292_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11293_/X
+ sky130_fd_sc_hd__o211a_1
X_13032_ _13056_/C _13030_/X _13039_/A vssd1 vssd1 vccd1 vccd1 _13032_/Y sky130_fd_sc_hd__o21ai_1
Xhold5370 _12043_/X vssd1 vssd1 vccd1 vccd1 _17171_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10244_ hold2499/X _16572_/Q _10610_/C vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__mux2_1
Xhold5381 _17049_/Q vssd1 vssd1 vccd1 vccd1 hold5381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5392 _10801_/X vssd1 vssd1 vccd1 vccd1 _16757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _17893_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4680 _16888_/Q vssd1 vssd1 vccd1 vccd1 hold4680/X sky130_fd_sc_hd__dlygate4sd3_1
X_10175_ hold2882/X hold4777/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__mux2_1
Xhold4691 _11554_/X vssd1 vssd1 vccd1 vccd1 _17008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3990 _15243_/X vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17771_ _17900_/CLK hold246/X vssd1 vssd1 vccd1 vccd1 _17771_/Q sky130_fd_sc_hd__dfxtp_1
X_14983_ hold1595/X _15006_/B _14982_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _14983_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout180 _11171_/B vssd1 vssd1 vccd1 vccd1 _11735_/B sky130_fd_sc_hd__buf_4
Xfanout191 _13886_/B vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__buf_4
X_16722_ _18053_/CLK _16722_/D vssd1 vssd1 vccd1 vccd1 _16722_/Q sky130_fd_sc_hd__dfxtp_1
X_13934_ hold730/X _17775_/Q _13942_/S vssd1 vssd1 vccd1 vccd1 hold731/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _18266_/CLK _16653_/D vssd1 vssd1 vccd1 vccd1 _16653_/Q sky130_fd_sc_hd__dfxtp_1
X_13865_ _17742_/Q _13868_/B _13865_/C vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _17252_/CLK _15604_/D vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _12825_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _17448_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16584_ _18235_/CLK _16584_/D vssd1 vssd1 vccd1 vccd1 _16584_/Q sky130_fd_sc_hd__dfxtp_1
X_13796_ hold2814/X hold4089/X _13796_/S vssd1 vssd1 vccd1 vccd1 _13797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ _18324_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _15535_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12747_ _12753_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _17425_/D sky130_fd_sc_hd__and2_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18382_/CLK hold823/X vssd1 vssd1 vccd1 vccd1 hold822/A sky130_fd_sc_hd__dfxtp_1
X_15466_ _15960_/Q _09386_/A _09386_/D hold349/X vssd1 vssd1 vccd1 vccd1 _15471_/B
+ sky130_fd_sc_hd__a22o_1
X_12678_ _12876_/A _12678_/B vssd1 vssd1 vccd1 vccd1 _17402_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17205_ _17205_/CLK _17205_/D vssd1 vssd1 vccd1 vccd1 _17205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11629_ hold4355/X _11726_/B _11628_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11629_/X
+ sky130_fd_sc_hd__o211a_1
X_14417_ hold129/X _14445_/B vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18185_ _18185_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15397_ hold397/X _15479_/A2 _15484_/B1 hold434/X _15396_/X vssd1 vssd1 vccd1 vccd1
+ _15402_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17136_ _17908_/CLK _17136_/D vssd1 vssd1 vccd1 vccd1 _17136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14348_ _14388_/A _14348_/B vssd1 vssd1 vccd1 vccd1 _17973_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold606 hold606/A vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 hold617/A vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 input70/X vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 hold639/A vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ _17884_/CLK _17067_/D vssd1 vssd1 vccd1 vccd1 _17067_/Q sky130_fd_sc_hd__dfxtp_1
X_14279_ hold1870/X _14272_/B _14278_/X _14546_/C1 vssd1 vssd1 vccd1 vccd1 _14279_/X
+ sky130_fd_sc_hd__o211a_1
X_16018_ _17524_/CLK _16018_/D vssd1 vssd1 vccd1 vccd1 hold704/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ hold219/X hold595/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__mux2_1
Xhold2007 _08483_/X vssd1 vssd1 vccd1 vccd1 _15870_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2018 _16220_/Q vssd1 vssd1 vccd1 vccd1 hold2018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _08318_/X vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1306 _18011_/Q vssd1 vssd1 vccd1 vccd1 hold1306/X sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ hold5/X hold469/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__mux2_1
Xhold1317 _18389_/Q vssd1 vssd1 vccd1 vccd1 hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 _15849_/Q vssd1 vssd1 vccd1 vccd1 hold1328/X sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _18025_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1339 la_data_in[6] vssd1 vssd1 vccd1 vccd1 hold1339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09323_ _15545_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09323_/Y sky130_fd_sc_hd__nand2_1
X_09254_ _12813_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _16238_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ _15539_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08205_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09185_ hold2928/X _09218_/B _09184_/X _12777_/A vssd1 vssd1 vccd1 vccd1 _09185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08136_ hold265/X hold355/X hold196/X vssd1 vssd1 vccd1 vccd1 _08137_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08067_ hold2727/X _08082_/B _08066_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _08067_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3220 _10231_/X vssd1 vssd1 vccd1 vccd1 _16567_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3231 _11911_/X vssd1 vssd1 vccd1 vccd1 _17127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3242 _17164_/Q vssd1 vssd1 vccd1 vccd1 hold3242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3253 _17379_/Q vssd1 vssd1 vccd1 vccd1 hold3253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3264 _09742_/X vssd1 vssd1 vccd1 vccd1 _16404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2530 _16176_/Q vssd1 vssd1 vccd1 vccd1 hold2530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3275 _16785_/Q vssd1 vssd1 vccd1 vccd1 hold3275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2541 _16236_/Q vssd1 vssd1 vccd1 vccd1 hold2541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3286 _09850_/X vssd1 vssd1 vccd1 vccd1 _16440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2552 _14123_/X vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3297 _17360_/Q vssd1 vssd1 vccd1 vccd1 hold3297/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17981_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08969_ hold184/X hold722/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__mux2_1
Xhold2563 _08412_/X vssd1 vssd1 vccd1 vccd1 _15836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2574 _15674_/Q vssd1 vssd1 vccd1 vccd1 hold2574/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1840 _16195_/Q vssd1 vssd1 vccd1 vccd1 hold1840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2585 _14835_/X vssd1 vssd1 vccd1 vccd1 _18207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1851 _08267_/X vssd1 vssd1 vccd1 vccd1 _15768_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ hold4445/X _13871_/B _11979_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11980_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2596 _17972_/Q vssd1 vssd1 vccd1 vccd1 hold2596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1862 _07979_/X vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 _14231_/X vssd1 vssd1 vccd1 vccd1 _17917_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1884 _13016_/X vssd1 vssd1 vccd1 vccd1 _17516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1895 _09322_/X vssd1 vssd1 vccd1 vccd1 _16271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10931_ _18004_/Q hold4353/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13650_ _13764_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13650_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ hold1248/X _16778_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _16276_/Q _17378_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13581_ _13758_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__or2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ hold2740/X _16755_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__mux2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ hold310/X _15486_/A2 _15446_/B1 hold448/X vssd1 vssd1 vccd1 vccd1 _15320_/X
+ sky130_fd_sc_hd__a22o_1
X_12532_ hold1868/X _17355_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__mux2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ hold126/X _08598_/B _08999_/B _12462_/X _15491_/A vssd1 vssd1 vccd1 vccd1
+ hold127/A sky130_fd_sc_hd__o311a_1
X_15251_ _16289_/Q _15477_/A2 _15487_/B1 hold425/X _15250_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_152_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ hold1625/X _16962_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__mux2_1
X_14202_ _14774_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__nand2_1
X_15182_ _15182_/A hold656/X vssd1 vssd1 vccd1 vccd1 _15211_/B sky130_fd_sc_hd__or2_4
X_12394_ _15304_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _17290_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ hold1249/X _14148_/B _14132_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ hold2769/X hold4540/X _11732_/C vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14064_ _14511_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__or2_1
X_11276_ _17764_/Q hold5227/X _11762_/C vssd1 vssd1 vccd1 vccd1 _11277_/B sky130_fd_sc_hd__mux2_1
X_13015_ _15519_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__or2_1
X_10227_ _10521_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__or2_1
X_17823_ _17855_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_1
X_10158_ _10524_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17754_ _17754_/CLK _17754_/D vssd1 vssd1 vccd1 vccd1 _17754_/Q sky130_fd_sc_hd__dfxtp_1
X_14966_ _15508_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14966_/Y sky130_fd_sc_hd__nor2_2
X_10089_ _10563_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16705_ _18231_/CLK _16705_/D vssd1 vssd1 vccd1 vccd1 _16705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ _13917_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _17766_/D sky130_fd_sc_hd__and2_1
X_17685_ _17749_/CLK _17685_/D vssd1 vssd1 vccd1 vccd1 _17685_/Q sky130_fd_sc_hd__dfxtp_1
X_14897_ _14897_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__or2_2
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16636_ _18226_/CLK _16636_/D vssd1 vssd1 vccd1 vccd1 _16636_/Q sky130_fd_sc_hd__dfxtp_1
X_13848_ hold3196/X _13758_/A _13847_/X vssd1 vssd1 vccd1 vccd1 _13848_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16567_ _18221_/CLK _16567_/D vssd1 vssd1 vccd1 vccd1 _16567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13779_ _13779_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ _18339_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15518_ hold1313/X _15560_/A2 _15517_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _15518_/X
+ sky130_fd_sc_hd__o211a_1
X_16498_ _18373_/CLK _16498_/D vssd1 vssd1 vccd1 vccd1 _16498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _18339_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
X_15449_ hold330/X _15484_/A2 _15447_/X vssd1 vssd1 vccd1 vccd1 _15452_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18168_ _18226_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ _17279_/CLK _17119_/D vssd1 vssd1 vccd1 vccd1 _17119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold425 hold425/A vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _18131_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold436 hold463/X vssd1 vssd1 vccd1 vccd1 hold464/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 hold447/A vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ hold839/X _16471_/Q _10055_/C vssd1 vssd1 vccd1 vccd1 _09942_/B sky130_fd_sc_hd__mux2_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout905 hold783/X vssd1 vssd1 vccd1 vccd1 hold784/A sky130_fd_sc_hd__buf_6
Xfanout916 hold769/X vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__buf_4
Xfanout927 hold466/X vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__buf_8
X_09872_ hold1763/X hold3446/X _10628_/C vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 hold1097/X vssd1 vssd1 vccd1 vccd1 hold1098/A sky130_fd_sc_hd__buf_6
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _18262_/Q vssd1 vssd1 vccd1 vccd1 hold1103/X sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ _15334_/A hold444/X vssd1 vssd1 vccd1 vccd1 _16030_/D sky130_fd_sc_hd__and2_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 _15843_/Q vssd1 vssd1 vccd1 vccd1 hold1114/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _14496_/X vssd1 vssd1 vccd1 vccd1 _18045_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 _15643_/Q vssd1 vssd1 vccd1 vccd1 hold1136/X sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _15284_/A hold137/X vssd1 vssd1 vccd1 vccd1 _15997_/D sky130_fd_sc_hd__and2_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 _08499_/X vssd1 vssd1 vccd1 vccd1 _15878_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 hold1158/A vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__buf_8
Xhold1169 _17859_/Q vssd1 vssd1 vccd1 vccd1 hold1169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ hold53/X hold521/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__mux2_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_170_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18225_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09306_ hold2466/X _09338_/A2 _09305_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09306_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ _15513_/A hold3003/X _09277_/S vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _15551_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08119_ _08141_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09099_ hold1465/X _09106_/B _09098_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _09099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11130_ _11670_/A _11130_/B vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__or2_1
Xhold970 hold970/A vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__or2_1
Xhold3050 _17407_/Q vssd1 vssd1 vccd1 vccd1 hold3050/X sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ _11203_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10012_/Y sky130_fd_sc_hd__nor2_1
Xhold3061 _17501_/Q vssd1 vssd1 vccd1 vccd1 hold3061/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3072 _17387_/Q vssd1 vssd1 vccd1 vccd1 hold3072/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3083 _17451_/Q vssd1 vssd1 vccd1 vccd1 hold3083/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3094 _12650_/X vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2360 _14667_/X vssd1 vssd1 vccd1 vccd1 _18126_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14820_ _15213_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__or2_1
Xhold2371 _09308_/X vssd1 vssd1 vccd1 vccd1 _16264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2382 _15126_/X vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2393 _07985_/X vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 _18309_/Q vssd1 vssd1 vccd1 vccd1 hold1670/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ hold1403/X _14774_/B _14750_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14751_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1681 hold6028/X vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__buf_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ hold1930/X _17145_/Q _13388_/S vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__mux2_1
Xhold1692 hold6040/X vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__buf_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_258_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17731_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ hold4089/X _13814_/B _13701_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13702_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17470_ _17482_/CLK _17470_/D vssd1 vssd1 vccd1 vccd1 _17470_/Q sky130_fd_sc_hd__dfxtp_1
X_10914_ _11106_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__or2_1
X_14682_ _15129_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14682_/X sky130_fd_sc_hd__or2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ hold2243/X hold3740/X _13844_/C vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16421_ _18373_/CLK _16421_/D vssd1 vssd1 vccd1 vccd1 _16421_/Q sky130_fd_sc_hd__dfxtp_1
X_13633_ hold4325/X _13832_/B _13632_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13633_/X
+ sky130_fd_sc_hd__o211a_1
X_10845_ _11640_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ _18330_/CLK _16352_/D vssd1 vssd1 vccd1 vccd1 _16352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13564_ hold3560/X _13883_/B _13563_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13564_/X
+ sky130_fd_sc_hd__o211a_1
X_10776_ _11640_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15303_ _15490_/A1 _15295_/X _15302_/X _15490_/B1 hold4461/X vssd1 vssd1 vccd1 vccd1
+ _15303_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12515_ _07826_/A _12514_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__mux2_1
X_13495_ hold5136/X _13880_/B _13494_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16283_ _18462_/CLK _16283_/D vssd1 vssd1 vccd1 vccd1 _16283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _18054_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
X_12446_ _17316_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ hold2518/X _15221_/B _15233_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15234_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15165_ _15219_/A hold609/X vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__nand2_1
X_12377_ _17283_/Q _12377_/B _12377_/C vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _12018_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__or2_1
X_14116_ _14850_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__or2_1
X_15096_ hold937/X _15109_/B _15095_/X _15030_/A vssd1 vssd1 vccd1 vccd1 hold938/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14047_ hold1941/X _14036_/B _14046_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14047_/X
+ sky130_fd_sc_hd__o211a_1
X_11259_ _11652_/A _11259_/B vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _17901_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15998_ _17331_/CLK _15998_/D vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__dfxtp_1
X_17737_ _17737_/CLK _17737_/D vssd1 vssd1 vccd1 vccd1 _17737_/Q sky130_fd_sc_hd__dfxtp_1
X_14949_ hold865/X _14952_/B _14948_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 hold866/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ hold747/X _08500_/B vssd1 vssd1 vccd1 vccd1 _08470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17668_ _17669_/CLK _17668_/D vssd1 vssd1 vccd1 vccd1 _17668_/Q sky130_fd_sc_hd__dfxtp_1
X_16619_ _18268_/CLK _16619_/D vssd1 vssd1 vccd1 vccd1 _16619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _17697_/CLK _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09022_ hold136/X hold525/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold526/A sky130_fd_sc_hd__mux2_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5903 _16930_/Q vssd1 vssd1 vccd1 vccd1 hold5903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5914 _17549_/Q vssd1 vssd1 vccd1 vccd1 hold5914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 data_in[16] vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5925 _17532_/Q vssd1 vssd1 vccd1 vccd1 hold5925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5936 _17753_/Q vssd1 vssd1 vccd1 vccd1 hold5936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5947 hold6009/X vssd1 vssd1 vccd1 vccd1 hold5947/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5958 _18376_/Q vssd1 vssd1 vccd1 vccd1 hold5958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold85/X vssd1 vssd1 vccd1 vccd1 input45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__buf_8
Xhold255 input32/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5969 _18043_/Q vssd1 vssd1 vccd1 vccd1 hold5969/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _09924_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__or2_1
Xfanout702 _08887_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 _14362_/A vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout724 _08585_/A vssd1 vssd1 vccd1 vccd1 _14905_/C1 sky130_fd_sc_hd__buf_4
Xfanout735 _15050_/A vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout746 _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__buf_4
X_09855_ _09975_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__or2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 _14065_/C1 vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__buf_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _12256_/C1 vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__buf_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 _14191_/C1 vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ hold68/X hold644/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _10506_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__or2_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ hold35/X hold508/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__mux2_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 fanout337/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 hold730/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _12420_/A _08668_/B vssd1 vssd1 vccd1 vccd1 _15955_/D sky130_fd_sc_hd__and2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ hold23/X hold435/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__mux2_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10630_ _11218_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _10630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ hold3431/X _10568_/B _10560_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _10561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ hold3811/X _12204_/A _12299_/X vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__a21oi_1
X_13280_ _13273_/X _13279_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_17_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10492_ _10586_/A _10628_/B _10491_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _16654_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ _12243_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12162_ _13794_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11113_ hold5749/X _11789_/B _11112_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11113_/X
+ sky130_fd_sc_hd__o211a_1
X_12093_ _12093_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__or2_1
X_16970_ _17882_/CLK _16970_/D vssd1 vssd1 vccd1 vccd1 _16970_/Q sky130_fd_sc_hd__dfxtp_1
X_15921_ _18413_/CLK _15921_/D vssd1 vssd1 vccd1 vccd1 hold619/A sky130_fd_sc_hd__dfxtp_1
X_11044_ hold3477/X _11732_/B _11043_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _17647_/CLK _15852_/D vssd1 vssd1 vccd1 vccd1 _15852_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _08079_/X vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ hold1565/X _14822_/B _14802_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14803_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _17747_/CLK _15783_/D vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ hold3451/X _12994_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__mux2_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _17522_/CLK _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14735_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nor2_2
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11946_ _12234_/A _11946_/B vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__or2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17453_/CLK _17453_/D vssd1 vssd1 vccd1 vccd1 _17453_/Q sky130_fd_sc_hd__dfxtp_1
X_14665_ hold2248/X _14664_/B _14664_/Y _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14665_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _12267_/A _11877_/B vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__or2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16404_ _18382_/CLK _16404_/D vssd1 vssd1 vccd1 vccd1 _16404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ hold2028/X _17659_/Q _13808_/C vssd1 vssd1 vccd1 vccd1 _13617_/B sky130_fd_sc_hd__mux2_1
X_17384_ _18438_/CLK _17384_/D vssd1 vssd1 vccd1 vccd1 _17384_/Q sky130_fd_sc_hd__dfxtp_1
X_10828_ hold3991/X _11210_/B _10827_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10828_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14596_ _15205_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14596_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16335_ _18416_/CLK _16335_/D vssd1 vssd1 vccd1 vccd1 _16335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13547_ _15821_/Q hold4651/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__mux2_1
X_10759_ hold3892/X _11726_/B _10758_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _10759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16266_ _17496_/CLK _16266_/D vssd1 vssd1 vccd1 vccd1 _16266_/Q sky130_fd_sc_hd__dfxtp_1
X_13478_ hold2281/X hold4377/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18005_ _18032_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ _15217_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15217_/Y sky130_fd_sc_hd__nand2_1
X_12429_ hold251/X hold393/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__mux2_1
X_16197_ _17475_/CLK _16197_/D vssd1 vssd1 vccd1 vccd1 _16197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4509 _11395_/X vssd1 vssd1 vccd1 vccd1 _16955_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15148_ hold1246/X _15161_/B _15147_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15148_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3808 _17098_/Q vssd1 vssd1 vccd1 vccd1 hold3808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3819 _17117_/Q vssd1 vssd1 vccd1 vccd1 hold3819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07970_ _15539_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__or2_1
X_15079_ _15187_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09640_ hold5666/X _10016_/B _09639_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09640_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18304_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09571_ hold5040/X _10070_/B _09570_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09571_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08522_ _17518_/Q _13043_/C vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__nand2b_2
XFILLER_0_171_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ hold1208/X _08488_/B _08452_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ _14726_/A hold1842/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ _12426_/A hold675/X vssd1 vssd1 vccd1 vccd1 _16119_/D sky130_fd_sc_hd__and2_1
XFILLER_0_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5700 _09538_/X vssd1 vssd1 vccd1 vccd1 _16336_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5711 _16951_/Q vssd1 vssd1 vccd1 vccd1 hold5711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5722 _11575_/X vssd1 vssd1 vccd1 vccd1 _17015_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5733 _16797_/Q vssd1 vssd1 vccd1 vccd1 hold5733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5744 _11599_/X vssd1 vssd1 vccd1 vccd1 _17023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5755 hold5906/X vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__buf_1
Xhold5766 output84/X vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_12
Xhold5777 hold5916/X vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5788 output75/X vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_12
Xhold5799 hold5928/X vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout510 fanout523/X vssd1 vssd1 vccd1 vccd1 _10610_/C sky130_fd_sc_hd__clkbuf_4
Xfanout521 _10523_/S vssd1 vssd1 vccd1 vccd1 _10637_/C sky130_fd_sc_hd__clkbuf_8
X_09907_ hold3857/X _10001_/B _09906_/X _15050_/A vssd1 vssd1 vccd1 vccd1 _09907_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout532 _09218_/B vssd1 vssd1 vccd1 vccd1 _09216_/B sky130_fd_sc_hd__buf_4
Xfanout543 _08866_/S vssd1 vssd1 vccd1 vccd1 _08860_/S sky130_fd_sc_hd__buf_8
Xfanout554 _08283_/Y vssd1 vssd1 vccd1 vccd1 _08336_/A2 sky130_fd_sc_hd__buf_8
Xfanout565 _08048_/Y vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__clkbuf_8
Xfanout576 _07865_/B vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__clkbuf_8
Xfanout587 _13198_/B vssd1 vssd1 vccd1 vccd1 _13310_/B sky130_fd_sc_hd__clkbuf_8
X_09838_ hold5385/X _10028_/B _09837_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09838_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout598 _12589_/S vssd1 vssd1 vccd1 vccd1 _12910_/S sky130_fd_sc_hd__buf_4
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09769_ hold3388/X _10601_/B _09768_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09769_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12343_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _11800_/Y sky130_fd_sc_hd__nor2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12789_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _17436_/D sky130_fd_sc_hd__and2_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12301_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11731_/Y sky130_fd_sc_hd__nor2_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ hold2614/X _14487_/B _14449_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14450_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ hold5470/X _12338_/B _11661_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11662_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13401_ _13791_/A _13401_/B vssd1 vssd1 vccd1 vccd1 _13401_/X sky130_fd_sc_hd__or2_1
X_10613_ _10613_/A _10637_/B _10637_/C vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11593_ hold5361/X _11783_/B _11592_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11593_/X
+ sky130_fd_sc_hd__o211a_1
X_14381_ _15169_/A hold1938/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__mux2_1
X_16120_ _17343_/CLK _16120_/D vssd1 vssd1 vccd1 vccd1 hold476/A sky130_fd_sc_hd__dfxtp_1
X_10544_ hold764/X _16672_/Q _10640_/C vssd1 vssd1 vccd1 vccd1 _10545_/B sky130_fd_sc_hd__mux2_1
X_13332_ _13716_/A _13332_/B vssd1 vssd1 vccd1 vccd1 _13332_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ _18308_/CLK _16051_/D vssd1 vssd1 vccd1 vccd1 _16051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13263_ _13311_/A1 _13261_/X _13262_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13263_/X
+ sky130_fd_sc_hd__o211a_1
X_10475_ hold2584/X hold3502/X _10571_/C vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15002_ _15109_/A _15006_/B vssd1 vssd1 vccd1 vccd1 _15002_/Y sky130_fd_sc_hd__nand2_1
X_12214_ hold4643/X _12308_/B _12213_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12214_/X
+ sky130_fd_sc_hd__o211a_1
X_13194_ _17575_/Q _17109_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12145_ hold3368/X _12377_/B _12144_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17257_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12076_ hold4671/X _13871_/B _12075_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__o211a_1
X_16953_ _17894_/CLK _16953_/D vssd1 vssd1 vccd1 vccd1 _16953_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_273_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17870_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15904_ _17531_/CLK _15904_/D vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__dfxtp_1
X_11027_ _18036_/Q _16833_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _11028_/B sky130_fd_sc_hd__mux2_1
X_16884_ _18055_/CLK _16884_/D vssd1 vssd1 vccd1 vccd1 _16884_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_202_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18065_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _17686_/CLK _15835_/D vssd1 vssd1 vccd1 vccd1 _15835_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _17749_/CLK _15766_/D vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfxtp_1
X_12978_ _12987_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _17502_/D sky130_fd_sc_hd__and2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17506_/CLK _17505_/D vssd1 vssd1 vccd1 vccd1 _17505_/Q sky130_fd_sc_hd__dfxtp_1
X_14717_ hold2306/X _14720_/B _14716_/Y _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14717_/X
+ sky130_fd_sc_hd__o211a_1
X_11929_ hold3474/X _12311_/B _11928_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _11929_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15697_ _17900_/CLK _15697_/D vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17436_ _17439_/CLK _17436_/D vssd1 vssd1 vccd1 vccd1 _17436_/Q sky130_fd_sc_hd__dfxtp_1
X_14648_ _14988_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14648_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_28 _09494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17367_ _17494_/CLK _17367_/D vssd1 vssd1 vccd1 vccd1 _17367_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_39 _15221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ hold2691/X _14610_/B _14578_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16318_ _18460_/CLK _16318_/D vssd1 vssd1 vccd1 vccd1 _16318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17298_ _17300_/CLK _17298_/D vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5007 _17027_/Q vssd1 vssd1 vccd1 vccd1 hold5007/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16249_ _17691_/CLK _16249_/D vssd1 vssd1 vccd1 vccd1 _16249_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5018 _09664_/X vssd1 vssd1 vccd1 vccd1 _16378_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5029 _11827_/X vssd1 vssd1 vccd1 vccd1 _17099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput102 _13121_/A vssd1 vssd1 vccd1 vccd1 hold5813/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4306 _10255_/X vssd1 vssd1 vccd1 vccd1 _16575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xoutput113 hold5827/X vssd1 vssd1 vccd1 vccd1 hold5828/A sky130_fd_sc_hd__buf_6
Xhold4317 _16639_/Q vssd1 vssd1 vccd1 vccd1 hold4317/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput124 hold5873/X vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_12
Xhold4328 _10345_/X vssd1 vssd1 vccd1 vccd1 _16605_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput135 hold4461/X vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_12
Xoutput146 hold5881/X vssd1 vssd1 vccd1 vccd1 slv_enable sky130_fd_sc_hd__buf_12
Xhold4339 _17034_/Q vssd1 vssd1 vccd1 vccd1 hold4339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3605 _11166_/Y vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3616 _16714_/Q vssd1 vssd1 vccd1 vccd1 hold3616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3627 _10600_/Y vssd1 vssd1 vccd1 vccd1 _16690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3638 _11158_/Y vssd1 vssd1 vccd1 vccd1 _16876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2904 _14456_/X vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3649 _11178_/Y vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2915 _17942_/Q vssd1 vssd1 vccd1 vccd1 hold2915/X sky130_fd_sc_hd__dlygate4sd3_1
X_07953_ hold2836/X _07991_/A2 _07952_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07953_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2926 _18327_/Q vssd1 vssd1 vccd1 vccd1 hold2926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2937 _14241_/X vssd1 vssd1 vccd1 vccd1 _17921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2948 _14406_/X vssd1 vssd1 vccd1 vccd1 _18001_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2959 _18139_/Q vssd1 vssd1 vccd1 vccd1 hold2959/X sky130_fd_sc_hd__dlygate4sd3_1
X_07884_ hold816/X hold585/X vssd1 vssd1 vccd1 vccd1 _07884_/Y sky130_fd_sc_hd__nor2_1
X_09623_ hold2719/X hold3859/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__mux2_1
X_09554_ hold2787/X _13206_/A _10571_/C vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08505_ _14218_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09485_ hold1601/X hold5887/X _09484_/B vssd1 vssd1 vccd1 vccd1 _09485_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08436_ hold5974/X _08440_/A2 hold741/X _08383_/A vssd1 vssd1 vccd1 vccd1 hold742/A
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_77_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18421_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _15815_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ hold2811/X _08336_/A2 _08297_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _08298_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5530 _16422_/Q vssd1 vssd1 vccd1 vccd1 hold5530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5541 _11488_/X vssd1 vssd1 vccd1 vccd1 _16986_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10260_ _10548_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__or2_1
Xhold5552 _16490_/Q vssd1 vssd1 vccd1 vccd1 hold5552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5563 _09607_/X vssd1 vssd1 vccd1 vccd1 _16359_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5574 _16762_/Q vssd1 vssd1 vccd1 vccd1 hold5574/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4840 _16610_/Q vssd1 vssd1 vccd1 vccd1 hold4840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5585 _11002_/X vssd1 vssd1 vccd1 vccd1 _16824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4851 _13549_/X vssd1 vssd1 vccd1 vccd1 _17636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5596 _16760_/Q vssd1 vssd1 vccd1 vccd1 hold5596/X sky130_fd_sc_hd__dlygate4sd3_1
X_10191_ _10557_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4862 _17240_/Q vssd1 vssd1 vccd1 vccd1 hold4862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4873 _17670_/Q vssd1 vssd1 vccd1 vccd1 hold4873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4884 _10279_/X vssd1 vssd1 vccd1 vccd1 _16583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4895 _17178_/Q vssd1 vssd1 vccd1 vccd1 hold4895/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout340 _12443_/S vssd1 vssd1 vccd1 vccd1 _12439_/S sky130_fd_sc_hd__buf_8
Xfanout351 _08910_/S vssd1 vssd1 vccd1 vccd1 _08930_/S sky130_fd_sc_hd__buf_8
Xfanout362 _15507_/Y vssd1 vssd1 vccd1 vccd1 _15560_/A2 sky130_fd_sc_hd__buf_4
Xfanout373 hold301/X vssd1 vssd1 vccd1 vccd1 _15069_/S sky130_fd_sc_hd__clkbuf_8
X_13950_ hold892/X _13992_/B vssd1 vssd1 vccd1 vccd1 _13950_/X sky130_fd_sc_hd__or2_1
Xfanout384 _14822_/B vssd1 vssd1 vccd1 vccd1 _14828_/B sky130_fd_sc_hd__buf_6
Xfanout395 _14545_/B vssd1 vssd1 vccd1 vccd1 _14553_/B sky130_fd_sc_hd__clkbuf_8
X_12901_ hold1923/X _17478_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__mux2_1
X_13881_ hold3969/X _13791_/A _13880_/X vssd1 vssd1 vccd1 vccd1 _13881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _17205_/CLK _15620_/D vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ hold1511/X hold2340/X _12844_/S vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__or2_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ hold2710/X _17432_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__mux2_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15182_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14545_/B sky130_fd_sc_hd__or2_4
X_18270_ _18304_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ hold2344/X _17062_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11715_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15482_ _15482_/A _15482_/B vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__and2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12694_ hold982/X _17409_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__mux2_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17221_ _17221_/CLK _17221_/D vssd1 vssd1 vccd1 vccd1 _17221_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _15547_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14433_/Y sky130_fd_sc_hd__nand2_1
X_11645_ hold2762/X _17039_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17152_ _17216_/CLK _17152_/D vssd1 vssd1 vccd1 vccd1 _17152_/Q sky130_fd_sc_hd__dfxtp_1
Xinput15 hold74/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__buf_1
XFILLER_0_135_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14364_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _17981_/D sky130_fd_sc_hd__and2_1
Xinput26 input26/A vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
X_11576_ hold2666/X _17016_/Q _11672_/S vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
X_16103_ _18413_/CLK _16103_/D vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__dfxtp_1
Xinput48 input48/A vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_6
X_13315_ hold5025/X _12311_/B _13314_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _17558_/D
+ sky130_fd_sc_hd__o211a_1
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10527_ _10527_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17083_ _17908_/CLK _17083_/D vssd1 vssd1 vccd1 vccd1 _17083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14295_ hold689/X _14333_/A2 _14294_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 hold690/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ _17313_/CLK _16034_/D vssd1 vssd1 vccd1 vccd1 hold680/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13246_ _13246_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13246_/X sky130_fd_sc_hd__or2_1
X_10458_ _10527_/A _10458_/B vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13177_ _13177_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__and2_1
XFILLER_0_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10485_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ hold2689/X hold4985/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__mux2_1
X_17985_ _18337_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 hold911/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12059_ hold1484/X hold4877/X _13388_/S vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__mux2_1
X_16936_ _17879_/CLK _16936_/D vssd1 vssd1 vccd1 vccd1 _16936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16867_ _18070_/CLK _16867_/D vssd1 vssd1 vccd1 vccd1 _16867_/Q sky130_fd_sc_hd__dfxtp_1
X_15818_ _17697_/CLK hold124/X vssd1 vssd1 vccd1 vccd1 _15818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16798_ _18065_/CLK _16798_/D vssd1 vssd1 vccd1 vccd1 _16798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15749_ _17694_/CLK _15749_/D vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09270_ _09272_/A hold336/X vssd1 vssd1 vccd1 vccd1 hold337/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08221_ hold800/X _08225_/B vssd1 vssd1 vccd1 vccd1 _08221_/X sky130_fd_sc_hd__or2_1
X_17419_ _17419_/CLK _17419_/D vssd1 vssd1 vccd1 vccd1 _17419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ _18399_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _15557_/A hold2611/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08083_ hold2336/X _08088_/B _08082_/Y _13941_/A vssd1 vssd1 vccd1 vccd1 _08083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4103 _17070_/Q vssd1 vssd1 vccd1 vccd1 hold4103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4114 _11584_/X vssd1 vssd1 vccd1 vccd1 _17018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4125 _16623_/Q vssd1 vssd1 vccd1 vccd1 hold4125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_195_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18054_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4136 _13417_/X vssd1 vssd1 vccd1 vccd1 _17592_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4147 _16669_/Q vssd1 vssd1 vccd1 vccd1 hold4147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3402 _17723_/Q vssd1 vssd1 vccd1 vccd1 hold3402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3413 _17259_/Q vssd1 vssd1 vccd1 vccd1 _12305_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4158 _10399_/X vssd1 vssd1 vccd1 vccd1 _16623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_124_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18235_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4169 _17578_/Q vssd1 vssd1 vccd1 vccd1 hold4169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3424 _17507_/Q vssd1 vssd1 vccd1 vccd1 hold3424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3435 _17374_/Q vssd1 vssd1 vccd1 vccd1 hold3435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3446 _16448_/Q vssd1 vssd1 vccd1 vccd1 hold3446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2701 _16262_/Q vssd1 vssd1 vccd1 vccd1 hold2701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _14991_/X vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3457 _12998_/X vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08985_ hold50/X hold472/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08986_/B sky130_fd_sc_hd__mux2_1
Xhold2723 _17809_/Q vssd1 vssd1 vccd1 vccd1 hold2723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3468 _17420_/Q vssd1 vssd1 vccd1 vccd1 hold3468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2734 _18456_/Q vssd1 vssd1 vccd1 vccd1 hold2734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3479 _16838_/Q vssd1 vssd1 vccd1 vccd1 hold3479/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2745 _14719_/X vssd1 vssd1 vccd1 vccd1 _18151_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2756 _18396_/Q vssd1 vssd1 vccd1 vccd1 hold2756/X sky130_fd_sc_hd__dlygate4sd3_1
X_07936_ _15559_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07936_/X sky130_fd_sc_hd__or2_1
Xhold2767 _16200_/Q vssd1 vssd1 vccd1 vccd1 hold2767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2778 hold5801/X vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__clkbuf_4
Xhold2789 _15622_/Q vssd1 vssd1 vccd1 vccd1 hold2789/X sky130_fd_sc_hd__dlygate4sd3_1
X_07867_ _15545_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _09903_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__or2_1
X_07798_ _07804_/A _09342_/A _09339_/B hold2989/X vssd1 vssd1 vccd1 vccd1 _07798_/X
+ sky130_fd_sc_hd__o22a_1
X_09537_ _09987_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09472_/C _09472_/D _09472_/B vssd1 vssd1 vccd1 vccd1 _09470_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_164_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _15207_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08419_/X sky130_fd_sc_hd__or2_1
X_09399_ _15559_/A _14555_/C _09399_/C _09398_/X vssd1 vssd1 vccd1 vccd1 _09400_/C
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _12204_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _12093_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ hold4109/X _10643_/B _10311_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__o211a_1
X_13100_ hold3607/X _13099_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__mux2_1
X_11292_ _12051_/A _11292_/B vssd1 vssd1 vccd1 vccd1 _11292_/X sky130_fd_sc_hd__or2_1
X_14080_ _15533_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__or2_1
Xhold5360 _09757_/X vssd1 vssd1 vccd1 vccd1 _16409_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13031_ _13030_/X _13039_/A _13031_/C vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__and3b_1
Xhold5371 _16469_/Q vssd1 vssd1 vccd1 vccd1 hold5371/X sky130_fd_sc_hd__dlygate4sd3_1
X_10243_ hold4030/X _10643_/B _10242_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10243_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5382 _11581_/X vssd1 vssd1 vccd1 vccd1 _17017_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5393 _16896_/Q vssd1 vssd1 vccd1 vccd1 hold5393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4670 _12241_/X vssd1 vssd1 vccd1 vccd1 _17237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4681 _11098_/X vssd1 vssd1 vccd1 vccd1 _16856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10174_ hold4375/X _10558_/A2 _10173_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10174_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4692 _16386_/Q vssd1 vssd1 vccd1 vccd1 hold4692/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3980 _16355_/Q vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__dlygate4sd3_1
X_17770_ _17898_/CLK hold439/X vssd1 vssd1 vccd1 vccd1 _17770_/Q sky130_fd_sc_hd__dfxtp_1
X_14982_ _15197_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__or2_1
Xhold3991 _16798_/Q vssd1 vssd1 vccd1 vccd1 hold3991/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout170 _12314_/B vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__buf_4
Xfanout181 _11171_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__buf_4
Xfanout192 _13886_/B vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__buf_4
X_16721_ _18053_/CLK _16721_/D vssd1 vssd1 vccd1 vccd1 _16721_/Q sky130_fd_sc_hd__dfxtp_1
X_13933_ _13933_/A hold352/X vssd1 vssd1 vccd1 vccd1 _17774_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16652_ _18210_/CLK _16652_/D vssd1 vssd1 vccd1 vccd1 _16652_/Q sky130_fd_sc_hd__dfxtp_1
X_13864_ _13864_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _17283_/CLK _15603_/D vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ hold3113/X _12814_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__mux2_1
X_16583_ _18205_/CLK _16583_/D vssd1 vssd1 vccd1 vccd1 _16583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ hold4989/X _12311_/B _13794_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _17718_/D
+ sky130_fd_sc_hd__o211a_1
X_18322_ _18378_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ hold2407/X _15547_/B _15533_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _15534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ hold3033/X _12745_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18253_ _18389_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ hold227/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15465_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12677_ hold3016/X _12676_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ _17268_/CLK _17204_/D vssd1 vssd1 vccd1 vccd1 _17204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ hold2324/X hold209/X _14415_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18184_ _18216_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
X_11628_ _11631_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11628_/X sky130_fd_sc_hd__or2_1
X_15396_ _17343_/Q _09362_/C _09362_/D hold476/X vssd1 vssd1 vccd1 vccd1 _15396_/X
+ sky130_fd_sc_hd__a22o_1
X_17135_ _17263_/CLK _17135_/D vssd1 vssd1 vccd1 vccd1 _17135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ _15189_/A hold2920/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14348_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11559_ _11658_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 hold607/A vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__buf_4
Xhold618 hold618/A vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold629 hold629/A vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17066_ _17882_/CLK _17066_/D vssd1 vssd1 vccd1 vccd1 _17066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14726_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__or2_1
X_16017_ _18423_/CLK _16017_/D vssd1 vssd1 vccd1 vccd1 _16017_/Q sky130_fd_sc_hd__dfxtp_1
X_13229_ _13228_/X hold3754/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _15766_/Q vssd1 vssd1 vccd1 vccd1 hold2008/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _09217_/X vssd1 vssd1 vccd1 vccd1 _16220_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _14426_/X vssd1 vssd1 vccd1 vccd1 _18011_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08770_ _15364_/A hold76/X vssd1 vssd1 vccd1 vccd1 _16005_/D sky130_fd_sc_hd__and2_1
Xhold1318 _15214_/X vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _18025_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1329 _08438_/X vssd1 vssd1 vccd1 vccd1 _15849_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16919_ _17895_/CLK _16919_/D vssd1 vssd1 vccd1 vccd1 _16919_/Q sky130_fd_sc_hd__dfxtp_1
X_17899_ _17908_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ hold1894/X _09325_/B _09321_/Y _15506_/A vssd1 vssd1 vccd1 vccd1 _09322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ _15529_/A hold1898/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09254_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ hold2111/X _08209_/B _08203_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09184_ _15513_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_305_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17629_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08066_ _15525_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3210 _16557_/Q vssd1 vssd1 vccd1 vccd1 hold3210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3221 _16675_/Q vssd1 vssd1 vccd1 vccd1 hold3221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3232 _16816_/Q vssd1 vssd1 vccd1 vccd1 hold3232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3243 _11926_/X vssd1 vssd1 vccd1 vccd1 _17132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3254 _12608_/X vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2520 _16214_/Q vssd1 vssd1 vccd1 vccd1 hold2520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 _17484_/Q vssd1 vssd1 vccd1 vccd1 hold3265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2531 _09127_/X vssd1 vssd1 vccd1 vccd1 _16176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3276 _10789_/X vssd1 vssd1 vccd1 vccd1 _16753_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3287 _16412_/Q vssd1 vssd1 vccd1 vccd1 hold3287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2542 _16185_/Q vssd1 vssd1 vccd1 vccd1 hold2542/X sky130_fd_sc_hd__dlygate4sd3_1
X_08968_ _15454_/A _08968_/B vssd1 vssd1 vccd1 vccd1 _16101_/D sky130_fd_sc_hd__and2_1
Xhold2553 _15800_/Q vssd1 vssd1 vccd1 vccd1 hold2553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3298 _12551_/X vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2564 _17963_/Q vssd1 vssd1 vccd1 vccd1 hold2564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 _16219_/Q vssd1 vssd1 vccd1 vccd1 hold1830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2575 _08069_/X vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07919_ hold2010/X _07924_/B _07918_/Y _08153_/A vssd1 vssd1 vccd1 vccd1 _07919_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2586 _16182_/Q vssd1 vssd1 vccd1 vccd1 hold2586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1841 _09165_/X vssd1 vssd1 vccd1 vccd1 _16195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1852 _18101_/Q vssd1 vssd1 vccd1 vccd1 hold1852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 _17789_/Q vssd1 vssd1 vccd1 vccd1 hold2597/X sky130_fd_sc_hd__dlygate4sd3_1
X_08899_ _15374_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _16067_/D sky130_fd_sc_hd__and2_1
Xhold1863 _16248_/Q vssd1 vssd1 vccd1 vccd1 hold1863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1874 _17513_/Q vssd1 vssd1 vccd1 vccd1 hold1874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1885 _15583_/Q vssd1 vssd1 vccd1 vccd1 hold1885/X sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ hold5526/X _11216_/B _10929_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10930_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_92_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _16096_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold1896 _17853_/Q vssd1 vssd1 vccd1 vccd1 hold1896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17785_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10861_ hold5508/X _11156_/B _10860_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10861_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12600_ _12918_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _17376_/D sky130_fd_sc_hd__and2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ hold1275/X hold3552/X _13847_/C vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__mux2_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ hold5417/X _11210_/B _10791_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _10792_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12936_/A _12531_/B vssd1 vssd1 vccd1 vccd1 _17353_/D sky130_fd_sc_hd__and2_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ hold138/X _15486_/A2 _15446_/B1 _16054_/Q vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _17324_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12462_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ hold915/X _14202_/B _14200_/Y _13935_/A vssd1 vssd1 vccd1 vccd1 hold916/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11413_ hold4939/X _12341_/B _11412_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _15182_/A hold656/X vssd1 vssd1 vccd1 vccd1 _15181_/Y sky130_fd_sc_hd__nor2_2
X_12393_ hold26/X hold578/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__mux2_1
X_14132_ _14866_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14132_/X sky130_fd_sc_hd__or2_1
X_11344_ hold4425/X _11726_/B _11343_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _11344_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ hold1621/X _14105_/A2 _14062_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _14063_/X
+ sky130_fd_sc_hd__o211a_1
X_11275_ hold5604/X _11753_/B _11274_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11275_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5190 _09874_/X vssd1 vssd1 vccd1 vccd1 _16448_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13014_ hold1420/X _13003_/Y _13013_/X _12936_/A vssd1 vssd1 vccd1 vccd1 _13014_/X
+ sky130_fd_sc_hd__o211a_1
X_10226_ hold2342/X _16566_/Q _10646_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__mux2_1
X_10157_ hold1852/X hold3684/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__mux2_1
X_17822_ _18051_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ hold2439/X _14952_/B _14964_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__o211a_1
X_17753_ _17754_/CLK input71/X vssd1 vssd1 vccd1 vccd1 _17753_/Q sky130_fd_sc_hd__dfxtp_1
X_10088_ hold934/X hold3188/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__mux2_1
X_16704_ _18198_/CLK _16704_/D vssd1 vssd1 vccd1 vccd1 _16704_/Q sky130_fd_sc_hd__dfxtp_1
X_13916_ _15205_/A hold2877/X _13942_/S vssd1 vssd1 vccd1 vccd1 _13917_/B sky130_fd_sc_hd__mux2_1
X_17684_ _17748_/CLK _17684_/D vssd1 vssd1 vccd1 vccd1 _17684_/Q sky130_fd_sc_hd__dfxtp_1
X_14896_ _14897_/A hold656/X vssd1 vssd1 vccd1 vccd1 hold657/A sky130_fd_sc_hd__nor2_2
X_16635_ _18225_/CLK _16635_/D vssd1 vssd1 vccd1 vccd1 _16635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ _17736_/Q _13847_/B _13847_/C vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16566_ _18140_/CLK _16566_/D vssd1 vssd1 vccd1 vccd1 _16566_/Q sky130_fd_sc_hd__dfxtp_1
X_13778_ hold2085/X hold3564/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13779_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15517_ _15517_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__or2_1
X_18305_ _18305_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ _12813_/A _12729_/B vssd1 vssd1 vccd1 vccd1 _17419_/D sky130_fd_sc_hd__and2_1
X_16497_ _18378_/CLK _16497_/D vssd1 vssd1 vccd1 vccd1 _16497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18236_ _18236_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
X_15448_ hold415/X _15486_/A2 _15486_/B1 hold324/X vssd1 vssd1 vccd1 vccd1 _15448_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _18231_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ _15979_/Q _09365_/B _09392_/C hold190/X _15378_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 hold404/A vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ _17584_/CLK _17118_/D vssd1 vssd1 vccd1 vccd1 _17118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ _18206_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
Xhold426 hold426/A vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold437 hold465/X vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__buf_6
XFILLER_0_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17049_ _17769_/CLK _17049_/D vssd1 vssd1 vccd1 vccd1 _17049_/Q sky130_fd_sc_hd__dfxtp_1
X_09940_ hold5670/X _10016_/B _09939_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout906 _15123_/A vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__clkbuf_16
X_09871_ hold5048/X _10601_/B _09870_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09871_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 hold573/X vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__buf_8
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 hold466/X vssd1 vssd1 vccd1 vccd1 _15105_/A sky130_fd_sc_hd__clkbuf_16
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 hold129/X vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__buf_8
X_08822_ hold443/X _16030_/Q _08860_/S vssd1 vssd1 vccd1 vccd1 hold444/A sky130_fd_sc_hd__mux2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 _14951_/X vssd1 vssd1 vccd1 vccd1 _18262_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _08426_/X vssd1 vssd1 vccd1 vccd1 _15843_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _15588_/Q vssd1 vssd1 vccd1 vccd1 hold1126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _08004_/X vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ hold136/X _15997_/Q _08787_/S vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__mux2_1
Xhold1148 la_data_in[8] vssd1 vssd1 vccd1 vccd1 hold1148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _15033_/X vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _12422_/A _08684_/B vssd1 vssd1 vccd1 vccd1 _15963_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09305_ _14986_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ _12789_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _16229_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09167_ hold1917/X _09164_/B _09166_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _14517_/A hold1025/X hold196/X vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _15105_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08049_ hold816/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__or2_4
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 hold971/A vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ hold895/X _16844_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__mux2_1
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3040 hold5990/X vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__clkbuf_2
X_10011_ _13142_/A _09933_/A _10010_/X vssd1 vssd1 vccd1 vccd1 _10011_/Y sky130_fd_sc_hd__a21oi_1
Xhold3051 _12692_/X vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3062 _12974_/X vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3073 _17498_/Q vssd1 vssd1 vccd1 vccd1 hold3073/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3084 _17497_/Q vssd1 vssd1 vccd1 vccd1 hold3084/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3095 _17396_/Q vssd1 vssd1 vccd1 vccd1 hold3095/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2350 _18040_/Q vssd1 vssd1 vccd1 vccd1 hold2350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2361 _18019_/Q vssd1 vssd1 vccd1 vccd1 hold2361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2372 _18344_/Q vssd1 vssd1 vccd1 vccd1 hold2372/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 _15807_/Q vssd1 vssd1 vccd1 vccd1 hold2383/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _18062_/Q vssd1 vssd1 vccd1 vccd1 hold2394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1660 _14939_/X vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _15197_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__or2_1
Xhold1671 _18257_/Q vssd1 vssd1 vccd1 vccd1 hold1671/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1682 _09411_/X vssd1 vssd1 vccd1 vccd1 _16291_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ hold4639/X _11798_/B _11961_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1693 _09427_/X vssd1 vssd1 vccd1 vccd1 _16299_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13800_/A _13701_/B vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__or2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ hold2760/X hold4119/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__mux2_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14681_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14724_/B sky130_fd_sc_hd__or2_4
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ hold4919/X _12377_/B _11892_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _18399_/CLK _16420_/D vssd1 vssd1 vccd1 vccd1 _16420_/Q sky130_fd_sc_hd__dfxtp_1
X_13632_ _13737_/A _13632_/B vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844_ _17975_/Q hold4145/X _11735_/C vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_298_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16351_ _18392_/CLK _16351_/D vssd1 vssd1 vccd1 vccd1 _16351_/Q sky130_fd_sc_hd__dfxtp_1
X_13563_ _13788_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ hold2715/X _16749_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _10776_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_227_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15302_ _15489_/A _15302_/B _15302_/C _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ hold1089/X _17349_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12514_/X sky130_fd_sc_hd__mux2_1
X_16282_ _18462_/CLK _16282_/D vssd1 vssd1 vccd1 vccd1 _16282_/Q sky130_fd_sc_hd__dfxtp_1
X_13494_ _13791_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18021_ _18053_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or2_1
X_12445_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_151_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ hold2098/X hold609/X _15163_/Y _15060_/A vssd1 vssd1 vccd1 vccd1 _15164_/X
+ sky130_fd_sc_hd__o211a_1
X_12376_ _13888_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12376_/Y sky130_fd_sc_hd__nor2_1
X_14115_ hold2676/X hold587/X _14114_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14115_/X
+ sky130_fd_sc_hd__o211a_1
X_11327_ hold2670/X hold4431/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__mux2_1
X_15095_ hold747/X _15125_/B vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _14726_/A _14050_/B vssd1 vssd1 vccd1 vccd1 _14046_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ hold2919/X hold3702/X _11747_/C vssd1 vssd1 vccd1 vccd1 _11259_/B sky130_fd_sc_hd__mux2_1
X_10209_ _10563_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11189_ _11189_/A _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__and3_1
X_17805_ _17891_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _17331_/CLK _15997_/D vssd1 vssd1 vccd1 vccd1 _15997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _15109_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nand2_1
X_17736_ _17736_/CLK _17736_/D vssd1 vssd1 vccd1 vccd1 _17736_/Q sky130_fd_sc_hd__dfxtp_1
X_17667_ _17731_/CLK _17667_/D vssd1 vssd1 vccd1 vccd1 _17667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14879_ hold855/X _14882_/B _14878_/Y _14879_/C1 vssd1 vssd1 vccd1 vccd1 hold856/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _18353_/CLK _16618_/D vssd1 vssd1 vccd1 vccd1 _16618_/Q sky130_fd_sc_hd__dfxtp_1
X_17598_ _17726_/CLK _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16549_ _18267_/CLK _16549_/D vssd1 vssd1 vccd1 vccd1 _16549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _16127_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18219_ _18219_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5904 _17528_/Q vssd1 vssd1 vccd1 vccd1 hold5904/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5915 _17531_/Q vssd1 vssd1 vccd1 vccd1 hold5915/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5926 _17541_/Q vssd1 vssd1 vccd1 vccd1 hold5926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold212 hold19/X vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5937 hold5993/X vssd1 vssd1 vccd1 vccd1 hold5937/X sky130_fd_sc_hd__buf_1
Xhold223 hold332/X vssd1 vssd1 vccd1 vccd1 hold333/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5948 _18248_/Q vssd1 vssd1 vccd1 vccd1 hold5948/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 input45/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5959 _18274_/Q vssd1 vssd1 vccd1 vccd1 hold5959/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold581/X vssd1 vssd1 vccd1 vccd1 hold582/A sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ hold1525/X _16465_/Q _10025_/C vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__mux2_1
Xhold289 hold37/X vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _09047_/A vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__clkbuf_4
Xfanout714 _14362_/A vssd1 vssd1 vccd1 vccd1 _14907_/C1 sky130_fd_sc_hd__buf_4
Xfanout725 _09063_/A vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__clkbuf_4
Xfanout736 _14985_/C1 vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__buf_4
X_09854_ hold1758/X hold3548/X _10271_/S vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__mux2_1
Xfanout747 fanout763/X vssd1 vssd1 vccd1 vccd1 _13681_/C1 sky130_fd_sc_hd__buf_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout758 _14065_/C1 vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__buf_4
Xfanout769 _12256_/C1 vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__buf_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _15284_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _16021_/D sky130_fd_sc_hd__and2_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ hold937/X _16419_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _09786_/B sky130_fd_sc_hd__mux2_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _12420_/A hold494/X vssd1 vssd1 vccd1 vccd1 _15988_/D sky130_fd_sc_hd__and2_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 hold770/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ hold68/X hold550/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08668_/B sky130_fd_sc_hd__mux2_1
XANTENNA_129 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _12380_/A _08598_/B vssd1 vssd1 vccd1 vccd1 _08619_/S sky130_fd_sc_hd__or2_2
XFILLER_0_193_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_320_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _10560_/A _10560_/B vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09219_ hold1879/X _09218_/B _09218_/Y _12831_/A vssd1 vssd1 vccd1 vccd1 _09219_/X
+ sky130_fd_sc_hd__o211a_1
X_10491_ _10491_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__or2_1
X_12230_ hold2399/X hold4502/X _13871_/C vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ hold2260/X _17211_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _11694_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__or2_1
X_12092_ hold1251/X _17188_/Q _12320_/C vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__mux2_1
Xhold790 hold790/A vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
X_15920_ _17751_/CLK _15920_/D vssd1 vssd1 vccd1 vccd1 hold523/A sky130_fd_sc_hd__dfxtp_1
X_11043_ _11637_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__or2_1
X_15851_ _17678_/CLK _15851_/D vssd1 vssd1 vccd1 vccd1 _15851_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2180 _18195_/Q vssd1 vssd1 vccd1 vccd1 hold2180/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _15195_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__or2_1
Xhold2191 _18178_/Q vssd1 vssd1 vccd1 vccd1 hold2191/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782_ _17649_/CLK _15782_/D vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ hold2697/X _17509_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__mux2_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 _14793_/X vssd1 vssd1 vccd1 vccd1 _18186_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17521_ _17522_/CLK _17521_/D vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ hold2056/X _14720_/B _14732_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14733_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ hold2189/X hold5348/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17456_/CLK _17452_/D vssd1 vssd1 vccd1 vccd1 _17452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _15219_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__nand2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ hold369/X hold3897/X _12356_/C vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__mux2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _18386_/CLK _16403_/D vssd1 vssd1 vccd1 vccd1 _16403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ hold4333/X _13805_/B _13614_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13615_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17383_ _18441_/CLK _17383_/D vssd1 vssd1 vccd1 vccd1 _17383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ _11667_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__or2_1
X_14595_ hold1797/X _14610_/B _14594_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14595_/X
+ sky130_fd_sc_hd__o211a_1
X_16334_ _18424_/CLK _16334_/D vssd1 vssd1 vccd1 vccd1 _16334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13546_ hold4259/X _13832_/B _13545_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13546_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ _11631_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16265_ _17496_/CLK _16265_/D vssd1 vssd1 vccd1 vccd1 _16265_/Q sky130_fd_sc_hd__dfxtp_1
X_13477_ hold5195/X _13859_/B _13476_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _11652_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15216_ hold1004/X _15219_/B _15215_/Y _15216_/C1 vssd1 vssd1 vccd1 vccd1 _15216_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18004_ _18069_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
X_12428_ _12428_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _17307_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16196_ _17475_/CLK _16196_/D vssd1 vssd1 vccd1 vccd1 _16196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ hold883/X _15149_/B vssd1 vssd1 vccd1 vccd1 _15147_/X sky130_fd_sc_hd__or2_1
X_12359_ _17277_/Q _13871_/B _13871_/C vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3809 _12303_/Y vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__dlygate4sd3_1
X_15078_ hold1690/X _15113_/B _15077_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15078_/X
+ sky130_fd_sc_hd__o211a_1
X_14029_ hold1754/X _14040_/B _14028_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14029_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ _09951_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__or2_1
X_08521_ _08868_/B _13056_/C _17520_/Q vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__or3b_1
X_17719_ _17719_/CLK _17719_/D vssd1 vssd1 vccd1 vccd1 _17719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_149_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08452_ hold892/X _08500_/B vssd1 vssd1 vccd1 vccd1 _08452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _15823_/D sky130_fd_sc_hd__and2_1
XFILLER_0_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09004_ hold407/X hold674/X _09062_/S vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__mux2_1
Xhold5701 _16392_/Q vssd1 vssd1 vccd1 vccd1 hold5701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5712 _11287_/X vssd1 vssd1 vccd1 vccd1 _16919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5723 _16879_/Q vssd1 vssd1 vccd1 vccd1 hold5723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5734 _10825_/X vssd1 vssd1 vccd1 vccd1 _16765_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5745 _16470_/Q vssd1 vssd1 vccd1 vccd1 hold5745/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5756 output98/X vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_12
Xhold5767 hold5912/X vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5778 output76/X vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_12
Xhold5789 hold5923/X vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout500 fanout523/X vssd1 vssd1 vccd1 vccd1 _10562_/S sky130_fd_sc_hd__buf_4
Xfanout511 _10067_/C vssd1 vssd1 vccd1 vccd1 _10271_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09906_ _09948_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__or2_1
Xfanout522 fanout523/X vssd1 vssd1 vccd1 vccd1 _10523_/S sky130_fd_sc_hd__buf_4
Xfanout533 _09178_/Y vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__buf_4
Xfanout544 _08498_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__clkbuf_8
Xfanout555 _08260_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__clkbuf_8
Xfanout566 _08043_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__buf_6
X_09837_ _09918_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__or2_1
Xfanout577 _07829_/Y vssd1 vssd1 vccd1 vccd1 _07865_/B sky130_fd_sc_hd__buf_6
Xfanout588 _13230_/B vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__clkbuf_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 _12982_/S vssd1 vssd1 vccd1 vccd1 _12955_/S sky130_fd_sc_hd__clkbuf_8
X_09768_ _10098_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__or2_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ hold44/X hold312/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08720_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _11067_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__or2_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ hold3737/X _11637_/A _11729_/X vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _12051_/A _11661_/B vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__or2_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ hold1866/X hold3969/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ _11194_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__nor2_1
X_14380_ _14380_/A hold423/X vssd1 vssd1 vccd1 vccd1 _17989_/D sky130_fd_sc_hd__and2_1
X_11592_ _11688_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_181_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ hold1828/X hold3883/X _13811_/C vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ hold4209/X _10631_/B _10542_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16050_ _18414_/CLK _16050_/D vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ _13262_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13262_/X sky130_fd_sc_hd__or2_1
X_10474_ hold4832/X _10568_/B _10473_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15001_ hold2074/X _15004_/B _15000_/Y _15066_/A vssd1 vssd1 vccd1 vccd1 _15001_/X
+ sky130_fd_sc_hd__o211a_1
X_12213_ _13797_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__or2_1
X_13193_ _13193_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__and2_1
XFILLER_0_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12144_ _12282_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ _13392_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__or2_1
X_16952_ _17896_/CLK _16952_/D vssd1 vssd1 vccd1 vccd1 _16952_/Q sky130_fd_sc_hd__dfxtp_1
X_15903_ _16128_/CLK _15903_/D vssd1 vssd1 vccd1 vccd1 hold709/A sky130_fd_sc_hd__dfxtp_1
X_11026_ hold5520/X _11216_/B _11025_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _11026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ _18054_/CLK _16883_/D vssd1 vssd1 vccd1 vccd1 _16883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _17634_/CLK _15834_/D vssd1 vssd1 vccd1 vccd1 _15834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _17708_/CLK _15765_/D vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfxtp_1
X_12977_ hold3097/X _12976_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__mux2_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_242_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17748_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17506_/CLK _17504_/D vssd1 vssd1 vccd1 vccd1 _17504_/Q sky130_fd_sc_hd__dfxtp_1
X_14716_ _15217_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14716_/Y sky130_fd_sc_hd__nand2_1
X_11928_ _13794_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15696_ _17908_/CLK _15696_/D vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ hold2277/X _14664_/B _14646_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14647_/X
+ sky130_fd_sc_hd__o211a_1
X_17435_ _17435_/CLK _17435_/D vssd1 vssd1 vccd1 vccd1 _17435_/Q sky130_fd_sc_hd__dfxtp_1
X_11859_ _12051_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14578_ _14740_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_29 _09494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _17494_/CLK _17366_/D vssd1 vssd1 vccd1 vccd1 _17366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13529_ hold1633/X hold3422/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16317_ _18460_/CLK _16317_/D vssd1 vssd1 vccd1 vccd1 _16317_/Q sky130_fd_sc_hd__dfxtp_1
X_17297_ _18425_/CLK _17297_/D vssd1 vssd1 vccd1 vccd1 hold663/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16248_ _17691_/CLK _16248_/D vssd1 vssd1 vccd1 vccd1 _16248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5008 _11515_/X vssd1 vssd1 vccd1 vccd1 _16995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5019 _17242_/Q vssd1 vssd1 vccd1 vccd1 hold5019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput103 _13129_/A vssd1 vssd1 vccd1 vccd1 hold5784/A sky130_fd_sc_hd__buf_6
XFILLER_0_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput114 hold5854/X vssd1 vssd1 vccd1 vccd1 hold5855/A sky130_fd_sc_hd__buf_6
XFILLER_0_3_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16179_ _17464_/CLK _16179_/D vssd1 vssd1 vccd1 vccd1 _16179_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4307 _16382_/Q vssd1 vssd1 vccd1 vccd1 hold4307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4318 _10351_/X vssd1 vssd1 vccd1 vccd1 _16607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput125 hold5839/X vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_12
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput136 hold4867/X vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_12
Xhold4329 _16446_/Q vssd1 vssd1 vccd1 vccd1 hold4329/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3606 _11167_/Y vssd1 vssd1 vccd1 vccd1 _16879_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3617 _11151_/Y vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3628 _16535_/Q vssd1 vssd1 vccd1 vccd1 hold3628/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3639 _16539_/Q vssd1 vssd1 vccd1 vccd1 hold3639/X sky130_fd_sc_hd__clkbuf_2
Xhold2905 _18109_/Q vssd1 vssd1 vccd1 vccd1 hold2905/X sky130_fd_sc_hd__dlygate4sd3_1
X_07952_ _14246_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07952_/X sky130_fd_sc_hd__or2_1
Xhold2916 _14283_/X vssd1 vssd1 vccd1 vccd1 _17942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2927 _15086_/X vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2938 _18144_/Q vssd1 vssd1 vccd1 vccd1 hold2938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2949 _18002_/Q vssd1 vssd1 vccd1 vccd1 hold2949/X sky130_fd_sc_hd__dlygate4sd3_1
X_07883_ hold279/X hold606/A hold298/X hold624/A vssd1 vssd1 vccd1 vccd1 hold585/A
+ sky130_fd_sc_hd__or4bb_1
X_09622_ hold5454/X _10013_/B _09621_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__o211a_1
X_09553_ hold4522/X _10049_/B _09552_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _09553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08504_ _08504_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__or2_2
XFILLER_0_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ hold5887/X _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _16322_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_38_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08435_ hold730/X _08443_/B vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__or2_1
XFILLER_0_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08366_ _15535_/A hold1633/X hold122/X vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ _14246_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08297_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18462_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5520 _16864_/Q vssd1 vssd1 vccd1 vccd1 hold5520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5531 _09700_/X vssd1 vssd1 vccd1 vccd1 _16390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5542 _16458_/Q vssd1 vssd1 vccd1 vccd1 hold5542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5553 _09904_/X vssd1 vssd1 vccd1 vccd1 _16458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5564 _17206_/Q vssd1 vssd1 vccd1 vccd1 hold5564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4830 _16552_/Q vssd1 vssd1 vccd1 vccd1 hold4830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5575 _10720_/X vssd1 vssd1 vccd1 vccd1 _16730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4841 _10264_/X vssd1 vssd1 vccd1 vccd1 _16578_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ hold3105/X _16554_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__mux2_1
Xhold5586 _16748_/Q vssd1 vssd1 vccd1 vccd1 hold5586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4852 _16902_/Q vssd1 vssd1 vccd1 vccd1 hold4852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5597 _10714_/X vssd1 vssd1 vccd1 vccd1 _16728_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4863 _12154_/X vssd1 vssd1 vccd1 vccd1 _17208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4874 _13555_/X vssd1 vssd1 vccd1 vccd1 _17638_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4885 _16503_/Q vssd1 vssd1 vccd1 vccd1 hold4885/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout330 fanout337/X vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__buf_4
Xhold4896 _11968_/X vssd1 vssd1 vccd1 vccd1 _17146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout341 _12425_/S vssd1 vssd1 vccd1 vccd1 _12443_/S sky130_fd_sc_hd__buf_8
Xfanout352 _08730_/X vssd1 vssd1 vccd1 vccd1 _08787_/S sky130_fd_sc_hd__buf_8
Xfanout363 _15211_/B vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__clkbuf_8
Xfanout374 _15012_/B vssd1 vssd1 vccd1 vccd1 _15018_/B sky130_fd_sc_hd__clkbuf_8
Xfanout385 _14788_/Y vssd1 vssd1 vccd1 vccd1 _14822_/B sky130_fd_sc_hd__buf_8
Xfanout396 _14554_/A2 vssd1 vssd1 vccd1 vccd1 _14541_/B sky130_fd_sc_hd__buf_6
X_12900_ _14360_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _17476_/D sky130_fd_sc_hd__and2_1
X_13880_ _17747_/Q _13880_/B _13880_/C vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__and3_1
XFILLER_0_159_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12831_ _12831_/A _12831_/B vssd1 vssd1 vccd1 vccd1 _17453_/D sky130_fd_sc_hd__and2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ hold1854/X _15547_/B _15549_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _15550_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12813_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _17430_/D sky130_fd_sc_hd__and2_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _15182_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14501_/Y sky130_fd_sc_hd__nor2_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ hold4506/X _12305_/B _11712_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15481_ _15481_/A1 _15474_/X _15480_/X _15481_/B1 _18424_/Q vssd1 vssd1 vccd1 vccd1
+ _15481_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12693_ _12789_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _17407_/D sky130_fd_sc_hd__and2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17252_/CLK _17220_/D vssd1 vssd1 vccd1 vccd1 _17220_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ hold2660/X _14433_/B _14431_/Y _14907_/C1 vssd1 vssd1 vccd1 vccd1 _14432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ hold4103/X _11747_/B _11643_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _11644_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17151_ _17282_/CLK _17151_/D vssd1 vssd1 vccd1 vccd1 _17151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14363_ _15531_/A hold1248/X hold275/X vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__mux2_1
Xinput16 input16/A vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_11575_ hold5721/X _11765_/B _11574_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__o211a_1
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
X_16102_ _17528_/CLK _16102_/D vssd1 vssd1 vccd1 vccd1 hold722/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ _13794_/A _13314_/B vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__or2_1
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10526_ hold1559/X hold3305/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__mux2_1
Xinput49 input49/A vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
X_17082_ _17898_/CLK _17082_/D vssd1 vssd1 vccd1 vccd1 _17082_/Q sky130_fd_sc_hd__dfxtp_1
X_14294_ hold667/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _17331_/CLK _16033_/D vssd1 vssd1 vccd1 vccd1 _16033_/Q sky130_fd_sc_hd__dfxtp_1
X_13245_ _13244_/X hold3639/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__mux2_1
X_10457_ hold2022/X _16643_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13176_ _13169_/X _13175_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17540_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_161_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10388_ hold2191/X _16620_/Q _10625_/C vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12127_ hold4785/X _12356_/B _12126_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12127_/X
+ sky130_fd_sc_hd__o211a_1
X_17984_ _17984_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12058_ hold4820/X _11798_/B _12057_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _12058_/X
+ sky130_fd_sc_hd__o211a_1
X_16935_ _17879_/CLK _16935_/D vssd1 vssd1 vccd1 vccd1 _16935_/Q sky130_fd_sc_hd__dfxtp_1
X_11009_ hold2738/X hold4186/X _11201_/C vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16866_ _18069_/CLK _16866_/D vssd1 vssd1 vccd1 vccd1 _16866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15817_ _17731_/CLK _15817_/D vssd1 vssd1 vccd1 vccd1 hold913/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797_ _18032_/CLK _16797_/D vssd1 vssd1 vccd1 vccd1 _16797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _17718_/CLK _15748_/D vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15679_ _17870_/CLK _15679_/D vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ hold1859/X _08213_/B _08219_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _08220_/X
+ sky130_fd_sc_hd__o211a_1
X_17418_ _17419_/CLK _17418_/D vssd1 vssd1 vccd1 vccd1 _17418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18398_ _18398_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _15714_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17349_ _17513_/CLK _17349_/D vssd1 vssd1 vccd1 vccd1 _17349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08082_ _15000_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4104 _11644_/X vssd1 vssd1 vccd1 vccd1 _17038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4115 _16855_/Q vssd1 vssd1 vccd1 vccd1 hold4115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4126 _10303_/X vssd1 vssd1 vccd1 vccd1 _16591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4137 _16977_/Q vssd1 vssd1 vccd1 vccd1 hold4137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4148 _10441_/X vssd1 vssd1 vccd1 vccd1 _16637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3403 _13714_/X vssd1 vssd1 vccd1 vccd1 _17691_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3414 _12211_/X vssd1 vssd1 vccd1 vccd1 _17227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4159 _16851_/Q vssd1 vssd1 vccd1 vccd1 hold4159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3425 _12992_/X vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3436 _17352_/Q vssd1 vssd1 vccd1 vccd1 hold3436/X sky130_fd_sc_hd__dlygate4sd3_1
X_08984_ _12438_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _16109_/D sky130_fd_sc_hd__and2_1
Xhold3447 _09778_/X vssd1 vssd1 vccd1 vccd1 _16416_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2702 _09304_/X vssd1 vssd1 vccd1 vccd1 _16262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3458 _17434_/Q vssd1 vssd1 vccd1 vccd1 hold3458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 _18057_/Q vssd1 vssd1 vccd1 vccd1 hold2713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3469 _17450_/Q vssd1 vssd1 vccd1 vccd1 hold3469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2724 _14007_/X vssd1 vssd1 vccd1 vccd1 _17809_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2735 _15556_/X vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07935_ hold2137/X _07924_/B _07934_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _07935_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2746 _18170_/Q vssd1 vssd1 vccd1 vccd1 hold2746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2757 _15228_/X vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_164_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18218_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2768 _09175_/X vssd1 vssd1 vccd1 vccd1 _16200_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2779 _13047_/X vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07866_ hold1966/X _07865_/B _07865_/Y _08139_/A vssd1 vssd1 vccd1 vccd1 _07866_/X
+ sky130_fd_sc_hd__o211a_1
X_09605_ hold2633/X _16359_/Q _09998_/C vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07797_ _18459_/Q _07788_/Y _18460_/Q hold2989/X _11155_/A vssd1 vssd1 vccd1 vccd1
+ _07797_/X sky130_fd_sc_hd__a221o_1
X_09536_ hold2983/X _13158_/A _10022_/C vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _09472_/C _09472_/D _09466_/Y vssd1 vssd1 vccd1 vccd1 _16316_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08418_ hold5953/X _08440_/A2 _08417_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08418_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ hold606/A hold298/A hold270/X vssd1 vssd1 vccd1 vccd1 _09398_/X sky130_fd_sc_hd__and3_1
XFILLER_0_163_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08349_ _08349_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ hold1165/X _16944_/Q _12320_/C vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__mux2_1
Xhold6040 _16317_/Q vssd1 vssd1 vccd1 vccd1 hold6040/X sky130_fd_sc_hd__dlygate4sd3_1
X_10311_ _10548_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _17769_/Q hold5236/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ _13030_/A _13034_/D hold901/X vssd1 vssd1 vccd1 vccd1 _13030_/X sky130_fd_sc_hd__and3_1
Xhold5350 _16437_/Q vssd1 vssd1 vccd1 vccd1 hold5350/X sky130_fd_sc_hd__dlygate4sd3_1
X_10242_ _10485_/A _10242_/B vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__or2_1
Xhold5361 _17053_/Q vssd1 vssd1 vccd1 vccd1 hold5361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5372 _09841_/X vssd1 vssd1 vccd1 vccd1 _16437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5383 _16497_/Q vssd1 vssd1 vccd1 vccd1 hold5383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5394 _11122_/X vssd1 vssd1 vccd1 vccd1 _16864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4660 _11050_/X vssd1 vssd1 vccd1 vccd1 _16840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4671 _17214_/Q vssd1 vssd1 vccd1 vccd1 hold4671/X sky130_fd_sc_hd__dlygate4sd3_1
X_10173_ _10557_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4682 _17728_/Q vssd1 vssd1 vccd1 vccd1 hold4682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4693 _09592_/X vssd1 vssd1 vccd1 vccd1 _16354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3970 _13881_/Y vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14981_ hold2838/X _15004_/B _14980_/X _15473_/A vssd1 vssd1 vccd1 vccd1 _14981_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3981 _10074_/Y vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout160 _13808_/B vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__buf_4
Xfanout171 _09494_/X vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__clkbuf_4
Xhold3992 _10828_/X vssd1 vssd1 vccd1 vccd1 _16766_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16720_ _18052_/CLK _16720_/D vssd1 vssd1 vccd1 vccd1 _16720_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout182 _10852_/A2 vssd1 vssd1 vccd1 vccd1 _11171_/B sky130_fd_sc_hd__clkbuf_4
Xfanout193 fanout209/X vssd1 vssd1 vccd1 vccd1 _13886_/B sky130_fd_sc_hd__buf_4
X_13932_ hold173/X hold351/X hold244/X vssd1 vssd1 vccd1 vccd1 hold352/A sky130_fd_sc_hd__mux2_1
X_16651_ _18268_/CLK _16651_/D vssd1 vssd1 vccd1 vccd1 _16651_/Q sky130_fd_sc_hd__dfxtp_1
X_13863_ hold3138/X _13767_/A _13862_/X vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__a21oi_1
X_12814_ hold1355/X _17449_/Q _12814_/S vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux2_1
X_15602_ _17703_/CLK _15602_/D vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfxtp_1
X_13794_ _13794_/A _13794_/B vssd1 vssd1 vccd1 vccd1 _13794_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16582_ _18118_/CLK _16582_/D vssd1 vssd1 vccd1 vccd1 _16582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ _18353_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
X_12745_ _16246_/Q hold3027/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__mux2_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _15533_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15533_/X sky130_fd_sc_hd__or2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18252_ _18378_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
X_15464_ _15482_/A _15464_/B vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__and2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12676_ hold1223/X _17403_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
X_17203_ _17865_/CLK _17203_/D vssd1 vssd1 vccd1 vccd1 _17203_/Q sky130_fd_sc_hd__dfxtp_1
X_14415_ _14988_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11627_ hold2421/X _17033_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__mux2_1
X_18183_ _18183_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
X_15395_ _15395_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17134_ _17262_/CLK _17134_/D vssd1 vssd1 vccd1 vccd1 _17134_/Q sky130_fd_sc_hd__dfxtp_1
X_14346_ _14350_/A _14346_/B vssd1 vssd1 vccd1 vccd1 _17972_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11558_ hold2054/X hold5460/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__mux2_1
Xhold608 hold608/A vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__clkbuf_2
X_10509_ _10527_/A _10509_/B vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__or2_1
X_17065_ _18431_/CLK _17065_/D vssd1 vssd1 vccd1 vccd1 _17065_/Q sky130_fd_sc_hd__dfxtp_1
Xhold619 hold619/A vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ hold1475/X _14272_/B _14276_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14277_/X
+ sky130_fd_sc_hd__o211a_1
X_11489_ hold2975/X _16987_/Q _12320_/C vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__mux2_1
X_16016_ _17302_/CLK _16016_/D vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13228_ hold5263/X _13227_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13183_/A1 _13157_/X _13158_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13159_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 _08263_/X vssd1 vssd1 vccd1 vccd1 _15766_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _15712_/Q vssd1 vssd1 vccd1 vccd1 hold1308/X sky130_fd_sc_hd__dlygate4sd3_1
X_17967_ _18033_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1319 _17767_/Q vssd1 vssd1 vccd1 vccd1 hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16918_ _18064_/CLK _16918_/D vssd1 vssd1 vccd1 vccd1 _16918_/Q sky130_fd_sc_hd__dfxtp_1
X_17898_ _17898_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_16849_ _18020_/CLK _16849_/D vssd1 vssd1 vccd1 vccd1 _16849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _15543_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09252_ _12813_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _16237_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08203_ _15537_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ hold1101/X _09218_/B _09182_/X _12777_/A vssd1 vssd1 vccd1 vccd1 _09183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ _15539_/A hold1193/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08134_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ hold5955/X _08082_/B _08064_/X _08159_/A vssd1 vssd1 vccd1 vccd1 hold968/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3200 _12854_/X vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3211 _10105_/X vssd1 vssd1 vccd1 vccd1 _16525_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3222 _10459_/X vssd1 vssd1 vccd1 vccd1 _16643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3233 _10882_/X vssd1 vssd1 vccd1 vccd1 _16784_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3244 _17362_/Q vssd1 vssd1 vccd1 vccd1 hold3244/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3255 _17720_/Q vssd1 vssd1 vccd1 vccd1 hold3255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2510 _14081_/X vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2521 _09205_/X vssd1 vssd1 vccd1 vccd1 _16214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3266 _12923_/X vssd1 vssd1 vccd1 vccd1 _12924_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08967_ hold214/X hold620/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08968_/B sky130_fd_sc_hd__mux2_1
Xhold2532 _18292_/Q vssd1 vssd1 vccd1 vccd1 hold2532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3277 _17741_/Q vssd1 vssd1 vccd1 vccd1 hold3277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3288 _09670_/X vssd1 vssd1 vccd1 vccd1 _16380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2543 _09145_/X vssd1 vssd1 vccd1 vccd1 _16185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 _08334_/X vssd1 vssd1 vccd1 vccd1 _15800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3299 _16849_/Q vssd1 vssd1 vccd1 vccd1 hold3299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1820 _15795_/Q vssd1 vssd1 vccd1 vccd1 hold1820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 _14327_/X vssd1 vssd1 vccd1 vccd1 _17963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1831 _09215_/X vssd1 vssd1 vccd1 vccd1 _16219_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07918_ _15000_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07918_/Y sky130_fd_sc_hd__nand2_1
Xhold2576 _18322_/Q vssd1 vssd1 vccd1 vccd1 hold2576/X sky130_fd_sc_hd__dlygate4sd3_1
X_08898_ hold71/X hold647/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__mux2_1
Xhold1842 _15824_/Q vssd1 vssd1 vccd1 vccd1 hold1842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2587 _09139_/X vssd1 vssd1 vccd1 vccd1 _16182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 _14615_/X vssd1 vssd1 vccd1 vccd1 _18101_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 _13965_/X vssd1 vssd1 vccd1 vccd1 _17789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 _15838_/Q vssd1 vssd1 vccd1 vccd1 hold1864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1875 _13010_/X vssd1 vssd1 vccd1 vccd1 _17513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1886 _07876_/X vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07849_ _15527_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__or2_1
Xhold1897 _14097_/X vssd1 vssd1 vccd1 vccd1 _17853_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _11136_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _09903_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ _11115_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10791_/X sky130_fd_sc_hd__or2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ hold3481/X _12529_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__mux2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ hold47/X _12509_/A2 _12505_/A3 _12460_/X _09063_/A vssd1 vssd1 vccd1 vccd1
+ hold48/A sky130_fd_sc_hd__o311a_1
X_14200_ _14950_/A _14202_/B vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__nand2_1
X_11412_ _12246_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__or2_1
X_15180_ hold2459/X hold609/X _15179_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _15180_/X
+ sky130_fd_sc_hd__o211a_1
X_12392_ _12428_/A _12392_/B vssd1 vssd1 vccd1 vccd1 _17289_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ hold5973/X hold587/X hold748/X _13931_/A vssd1 vssd1 vccd1 vccd1 hold749/A
+ sky130_fd_sc_hd__o211a_1
X_11343_ _11631_/A _11343_/B vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _14850_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14062_/X sky130_fd_sc_hd__or2_1
X_11274_ _11658_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11274_/X sky130_fd_sc_hd__or2_1
Xhold5180 _13471_/X vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13013_ _15517_/A _13017_/B vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__or2_1
X_10225_ hold4073/X _10640_/B _10224_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10225_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5191 _16015_/Q vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4490 _17247_/Q vssd1 vssd1 vccd1 vccd1 hold4490/X sky130_fd_sc_hd__dlygate4sd3_1
X_17821_ _17856_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_1
X_10156_ hold4273/X _10646_/B _10155_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10156_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_4
X_17752_ _18462_/CLK _17752_/D vssd1 vssd1 vccd1 vccd1 _17752_/Q sky130_fd_sc_hd__dfxtp_1
X_10087_ hold5094/X _10568_/B _10086_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10087_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14964_ _15233_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_1
X_16703_ _18197_/CLK _16703_/D vssd1 vssd1 vccd1 vccd1 _16703_/Q sky130_fd_sc_hd__dfxtp_1
X_13915_ _14350_/A hold753/X vssd1 vssd1 vccd1 vccd1 _17765_/D sky130_fd_sc_hd__and2_1
X_17683_ _17737_/CLK _17683_/D vssd1 vssd1 vccd1 vccd1 _17683_/Q sky130_fd_sc_hd__dfxtp_1
X_14895_ hold2703/X _14882_/B _14894_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14895_/X
+ sky130_fd_sc_hd__o211a_1
X_16634_ _18192_/CLK _16634_/D vssd1 vssd1 vccd1 vccd1 _16634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ _13888_/A _13846_/B vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16565_ _18233_/CLK _16565_/D vssd1 vssd1 vccd1 vccd1 _16565_/Q sky130_fd_sc_hd__dfxtp_1
X_13777_ hold4747/X _13871_/B _13776_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__o211a_1
X_10989_ _11097_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10989_/X sky130_fd_sc_hd__or2_1
X_18304_ _18304_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ hold1529/X _15560_/A2 _15515_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _15516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ hold3486/X _12727_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _18399_/CLK _16496_/D vssd1 vssd1 vccd1 vccd1 _16496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18235_ _18235_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
X_15447_ hold725/X _15487_/B1 _15447_/B1 hold695/X vssd1 vssd1 vccd1 vccd1 _15447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ hold3095/X _12658_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ _18210_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
X_15378_ hold699/X _09386_/A _09392_/D hold353/X vssd1 vssd1 vccd1 vccd1 _15378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17117_ _17744_/CLK _17117_/D vssd1 vssd1 vccd1 vccd1 _17117_/Q sky130_fd_sc_hd__dfxtp_1
Xhold405 hold77/X vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14329_ hold2298/X _14333_/A2 _14328_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14329_/X
+ sky130_fd_sc_hd__o211a_1
Xhold416 hold416/A vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ _18225_/CLK hold940/X vssd1 vssd1 vccd1 vccd1 hold939/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold438 hold438/A vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _17896_/CLK _17048_/D vssd1 vssd1 vccd1 vccd1 _17048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09870_ _10506_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout907 _15123_/A vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__clkbuf_16
Xfanout918 hold573/X vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__buf_8
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 hold466/X vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__buf_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _12430_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _16029_/D sky130_fd_sc_hd__and2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 _15650_/Q vssd1 vssd1 vccd1 vccd1 hold1105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _17892_/Q vssd1 vssd1 vccd1 vccd1 hold1116/X sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _15344_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _15996_/D sky130_fd_sc_hd__and2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _07889_/X vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 _17886_/Q vssd1 vssd1 vccd1 vccd1 hold1138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 hold1149/A vssd1 vssd1 vccd1 vccd1 input67/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08683_ hold443/X hold672/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08684_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09304_ hold2701/X _09338_/A2 _09303_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ hold892/X hold982/X _09277_/S vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _15549_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08117_ _13929_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ hold2582/X _09106_/B _09096_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08048_ hold816/X _14627_/A vssd1 vssd1 vccd1 vccd1 _08048_/Y sky130_fd_sc_hd__nor2_2
Xhold950 hold950/A vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3030 _14693_/X vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _16494_/Q _10013_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__and3_1
Xhold3041 _12515_/X vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3052 _17439_/Q vssd1 vssd1 vccd1 vccd1 hold3052/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3063 _17458_/Q vssd1 vssd1 vccd1 vccd1 hold3063/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3074 _17384_/Q vssd1 vssd1 vccd1 vccd1 hold3074/X sky130_fd_sc_hd__dlygate4sd3_1
X_09999_ _13110_/A _09903_/A _09998_/X vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__a21oi_1
Xhold2340 _17455_/Q vssd1 vssd1 vccd1 vccd1 hold2340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3085 _17421_/Q vssd1 vssd1 vccd1 vccd1 hold3085/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3096 _12659_/X vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2351 _14486_/X vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2362 _14442_/X vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2373 _15120_/X vssd1 vssd1 vccd1 vccd1 _18344_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2384 _16224_/Q vssd1 vssd1 vccd1 vccd1 hold2384/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1650 _15763_/Q vssd1 vssd1 vccd1 vccd1 hold1650/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 _14532_/X vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ _12153_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__or2_1
Xhold1661 _17888_/Q vssd1 vssd1 vccd1 vccd1 hold1661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1672 _14941_/X vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1683 _17768_/Q vssd1 vssd1 vccd1 vccd1 hold1683/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 _15590_/Q vssd1 vssd1 vccd1 vccd1 hold1694/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ hold1850/X _17687_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13701_/B sky130_fd_sc_hd__mux2_1
X_10912_ hold5629/X _11213_/B _10911_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10912_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14681_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14680_/Y sky130_fd_sc_hd__nor2_1
X_11892_ _12282_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or2_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ hold1271/X hold4230/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__mux2_1
X_10843_ hold4248/X _11765_/B _10842_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _10843_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13562_ _15826_/Q hold3550/X _13886_/C vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _18385_/CLK _16350_/D vssd1 vssd1 vccd1 vccd1 _16350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ hold4045/X _11156_/B _10773_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _10774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15301_ _16294_/Q _15477_/A2 _15487_/B1 hold633/X _15300_/X vssd1 vssd1 vccd1 vccd1
+ _15302_/D sky130_fd_sc_hd__a221o_1
X_12513_ _13048_/A hold2175/X _07809_/X _18462_/Q vssd1 vssd1 vccd1 vccd1 _12513_/X
+ sky130_fd_sc_hd__a211o_1
X_16281_ _17751_/CLK _16281_/D vssd1 vssd1 vccd1 vccd1 _16281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ hold910/X hold5082/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18020_ _18020_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
X_12444_ _15284_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _17315_/D sky130_fd_sc_hd__and2_1
X_15232_ hold2957/X _15221_/B _15231_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_267_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _15217_/A hold609/X vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__nand2_1
X_12375_ hold3740/X _13749_/A _12374_/X vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _14740_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__or2_1
X_11326_ hold3392/X _11741_/B _11325_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__o211a_1
X_15094_ hold1486/X _15109_/B _15093_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15094_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14045_ hold1132/X _14036_/B _14044_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _14045_/X
+ sky130_fd_sc_hd__o211a_1
X_11257_ hold4369/X _11735_/B _11256_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ hold2880/X hold4657/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11188_ _11218_/A _11188_/B vssd1 vssd1 vccd1 vccd1 _11188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17804_ _17887_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_1
X_10139_ hold1844/X _16537_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__mux2_1
X_15996_ _18410_/CLK _15996_/D vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__dfxtp_1
X_17735_ _17735_/CLK _17735_/D vssd1 vssd1 vccd1 vccd1 _17735_/Q sky130_fd_sc_hd__dfxtp_1
X_14947_ hold1430/X _14946_/B _14946_/Y _15144_/C1 vssd1 vssd1 vccd1 vccd1 _14947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17666_ _17666_/CLK _17666_/D vssd1 vssd1 vccd1 vccd1 _17666_/Q sky130_fd_sc_hd__dfxtp_1
X_14878_ _15109_/A _14882_/B vssd1 vssd1 vccd1 vccd1 _14878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _18267_/CLK _16617_/D vssd1 vssd1 vccd1 vccd1 _16617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ _13829_/A _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__and3_1
X_17597_ _17629_/CLK _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _18228_/CLK _16548_/D vssd1 vssd1 vccd1 vccd1 _16548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _18392_/CLK _16479_/D vssd1 vssd1 vccd1 vccd1 _16479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ hold53/X hold327/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__mux2_1
X_18218_ _18218_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5905 _17527_/Q vssd1 vssd1 vccd1 vccd1 hold5905/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18149_ _18149_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5916 _17539_/Q vssd1 vssd1 vccd1 vccd1 hold5916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 hold34/X vssd1 vssd1 vccd1 vccd1 input30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5927 _17554_/Q vssd1 vssd1 vccd1 vccd1 hold5927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 input12/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5938 hold5995/X vssd1 vssd1 vccd1 vccd1 hold5938/X sky130_fd_sc_hd__buf_1
Xhold224 hold334/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__buf_6
Xhold5949 _17874_/Q vssd1 vssd1 vccd1 vccd1 hold5949/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold86/X vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__buf_4
XFILLER_0_1_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold279 hold583/X vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__clkbuf_8
X_09922_ hold5578/X _10016_/B _09921_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09922_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout704 _08887_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__clkbuf_4
Xfanout715 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__clkbuf_4
Xfanout726 _09063_/A vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__clkbuf_4
X_09853_ hold4047/X _10001_/B _09852_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09853_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout737 _08585_/A vssd1 vssd1 vccd1 vccd1 _14985_/C1 sky130_fd_sc_hd__buf_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08141_/A sky130_fd_sc_hd__buf_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 fanout763/X vssd1 vssd1 vccd1 vccd1 _14065_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ hold23/X hold324/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__mux2_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ hold4291/X _10070_/B _09783_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09784_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ hold407/X hold493/X _08793_/S vssd1 vssd1 vccd1 vccd1 hold494/A sky130_fd_sc_hd__mux2_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _14984_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _12428_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _15954_/D sky130_fd_sc_hd__and2_1
XANTENNA_119 hold770/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _17519_/Q _17518_/Q vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__nand2_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09218_ _15547_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ hold1499/X hold3204/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09149_ hold1130/X _09164_/B _09148_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _09149_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ hold5019/X _12347_/B _12159_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _12160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ hold2386/X hold4475/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__mux2_1
X_12091_ hold4486/X _12377_/B _12090_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12091_/X
+ sky130_fd_sc_hd__o211a_1
Xhold780 hold780/A vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold791 becStatus[3] vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ hold2155/X _16838_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__mux2_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _17741_/CLK _15850_/D vssd1 vssd1 vccd1 vccd1 _15850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2170 _17899_/Q vssd1 vssd1 vccd1 vccd1 hold2170/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2181 _14811_/X vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14801_ hold2995/X _14828_/B _14800_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14801_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _14775_/X vssd1 vssd1 vccd1 vccd1 _18178_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _17739_/CLK _15781_/D vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12996_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _17507_/D sky130_fd_sc_hd__and2_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _17522_/CLK _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1480 _18448_/Q vssd1 vssd1 vccd1 vccd1 hold1480/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1491 _17871_/Q vssd1 vssd1 vccd1 vccd1 hold1491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14732_ _14786_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__or2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ hold3495/X _13871_/B _11943_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17456_/CLK _17451_/D vssd1 vssd1 vccd1 vccd1 _17451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11875_ hold3521/X _12356_/B _11874_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _11875_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ hold2342/X _14666_/B _14662_/Y _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14663_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _18315_/CLK _16402_/D vssd1 vssd1 vccd1 vccd1 _16402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _13710_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13614_/X sky130_fd_sc_hd__or2_1
X_10826_ hold2096/X _16766_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _10827_/B sky130_fd_sc_hd__mux2_1
X_17382_ _18441_/CLK _17382_/D vssd1 vssd1 vccd1 vccd1 _17382_/Q sky130_fd_sc_hd__dfxtp_1
X_14594_ _14988_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14594_/X sky130_fd_sc_hd__or2_1
X_16333_ _18420_/CLK _16333_/D vssd1 vssd1 vccd1 vccd1 _16333_/Q sky130_fd_sc_hd__dfxtp_1
X_13545_ _13737_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__or2_1
X_10757_ hold2664/X _16743_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13476_ _13764_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _17494_/CLK _16264_/D vssd1 vssd1 vccd1 vccd1 _16264_/Q sky130_fd_sc_hd__dfxtp_1
X_10688_ hold2977/X hold3696/X _11747_/C vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__mux2_1
X_18003_ _18003_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
X_15215_ _15215_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15215_/Y sky130_fd_sc_hd__nand2_1
X_12427_ hold149/X hold191/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12428_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16195_ _17480_/CLK _16195_/D vssd1 vssd1 vccd1 vccd1 _16195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15146_ hold1286/X _15161_/B _15145_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _15146_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _13873_/A _12358_/B vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _17775_/Q hold5321/X _11789_/C vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__mux2_1
X_15077_ _15185_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__or2_1
X_12289_ hold4427/X _12308_/B _12288_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12289_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14028_ _15535_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15979_ _18414_/CLK _15979_/D vssd1 vssd1 vccd1 vccd1 _15979_/Q sky130_fd_sc_hd__dfxtp_1
X_08520_ _18460_/Q _13057_/B vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__nand2_1
X_17718_ _17718_/CLK _17718_/D vssd1 vssd1 vccd1 vccd1 _17718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ hold2781/X _08488_/B _08450_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08451_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17649_ _17649_/CLK _17649_/D vssd1 vssd1 vccd1 vccd1 _17649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08382_ _14330_/A hold1024/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_189_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18176_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_118_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18383_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _16118_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5702 _09610_/X vssd1 vssd1 vccd1 vccd1 _16360_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5713 _17087_/Q vssd1 vssd1 vccd1 vccd1 hold5713/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5724 _11071_/X vssd1 vssd1 vccd1 vccd1 _16847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5735 _16981_/Q vssd1 vssd1 vccd1 vccd1 hold5735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5746 _09844_/X vssd1 vssd1 vccd1 vccd1 _16438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5757 hold5907/X vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5768 output90/X vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_12
Xhold5779 hold5919/X vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout501 _10568_/C vssd1 vssd1 vccd1 vccd1 _10571_/C sky130_fd_sc_hd__clkbuf_8
X_09905_ hold2818/X hold3833/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__mux2_1
Xfanout512 _10067_/C vssd1 vssd1 vccd1 vccd1 _10628_/C sky130_fd_sc_hd__clkbuf_8
Xfanout523 _09499_/Y vssd1 vssd1 vccd1 vccd1 fanout523/X sky130_fd_sc_hd__clkbuf_8
Xfanout534 _09170_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__clkbuf_4
Xfanout545 _08448_/Y vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__clkbuf_8
Xfanout556 _08228_/Y vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__buf_8
X_09836_ hold1589/X hold3263/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__mux2_1
Xfanout567 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08029_/B sky130_fd_sc_hd__buf_8
Xfanout578 _14622_/B vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__clkbuf_8
Xfanout589 _13049_/Y vssd1 vssd1 vccd1 vccd1 _13183_/C1 sky130_fd_sc_hd__buf_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ hold1587/X _16413_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _15482_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _15980_/D sky130_fd_sc_hd__and2_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _18303_/Q hold5524/X _11066_/S vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__mux2_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ hold50/X hold168/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__mux2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ hold1116/X hold5367/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__mux2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ hold3135/X _10521_/A _10610_/X vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _17869_/Q hold5334/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__mux2_1
X_13330_ hold3396/X _13805_/B _13329_/X _12810_/A vssd1 vssd1 vccd1 vccd1 _13330_/X
+ sky130_fd_sc_hd__o211a_1
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13261_ _13260_/X hold3734/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _10560_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15000_ _15000_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15000_/Y sky130_fd_sc_hd__nand2_1
X_12212_ hold2388/X _17228_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _13185_/X _13191_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17542_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ hold2870/X _17205_/Q _12368_/C vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12074_ hold2516/X hold4445/X _13871_/C vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__mux2_1
X_16951_ _17895_/CLK _16951_/D vssd1 vssd1 vccd1 vccd1 _16951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15902_ _18421_/CLK _15902_/D vssd1 vssd1 vccd1 vccd1 hold557/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ _11121_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/X sky130_fd_sc_hd__or2_1
X_16882_ _18053_/CLK _16882_/D vssd1 vssd1 vccd1 vccd1 _16882_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _17724_/CLK _15833_/D vssd1 vssd1 vccd1 vccd1 _15833_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _17748_/CLK hold874/X vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__dfxtp_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ hold2048/X _17503_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__mux2_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17503_/CLK _17503_/D vssd1 vssd1 vccd1 vccd1 _17503_/Q sky130_fd_sc_hd__dfxtp_1
X_14715_ hold2070/X _14718_/B _14714_/Y _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14715_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ hold2727/X _17133_/Q _12353_/C vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__mux2_1
X_15695_ _17263_/CLK _15695_/D vssd1 vssd1 vccd1 vccd1 hold941/A sky130_fd_sc_hd__dfxtp_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17434_ _17435_/CLK _17434_/D vssd1 vssd1 vccd1 vccd1 _17434_/Q sky130_fd_sc_hd__dfxtp_1
X_14646_ _14986_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14646_/X sky130_fd_sc_hd__or2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ hold1203/X hold5278/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_282_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17856_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ _17494_/CLK _17365_/D vssd1 vssd1 vccd1 vccd1 _17365_/Q sky130_fd_sc_hd__dfxtp_1
X_10809_ _10998_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
X_14577_ hold1020/X _14612_/B _14576_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _14577_/X
+ sky130_fd_sc_hd__o211a_1
X_11789_ _17087_/Q _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__and3_1
XFILLER_0_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_211_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _17503_/CLK _16316_/D vssd1 vssd1 vccd1 vccd1 _16316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13528_ hold4417/X _13814_/B _13527_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _13528_/X
+ sky130_fd_sc_hd__o211a_1
X_17296_ _17318_/CLK _17296_/D vssd1 vssd1 vccd1 vccd1 hold698/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16247_ _17666_/CLK hold145/X vssd1 vssd1 vccd1 vccd1 _16247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ hold4826/X _13859_/B _13458_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13459_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5009 _16411_/Q vssd1 vssd1 vccd1 vccd1 hold5009/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput104 _10651_/A vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_12
Xoutput115 hold5874/X vssd1 vssd1 vccd1 vccd1 hold5875/A sky130_fd_sc_hd__buf_6
XFILLER_0_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16178_ _18441_/CLK _16178_/D vssd1 vssd1 vccd1 vccd1 _16178_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4308 _09580_/X vssd1 vssd1 vccd1 vccd1 _16350_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4319 _16424_/Q vssd1 vssd1 vccd1 vccd1 hold4319/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput126 hold5845/X vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_12
Xoutput137 hold5843/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_12
X_15129_ _15129_/A _15149_/B vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3607 _16713_/Q vssd1 vssd1 vccd1 vccd1 hold3607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3618 _11152_/Y vssd1 vssd1 vccd1 vccd1 _16874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3629 _10615_/Y vssd1 vssd1 vccd1 vccd1 _16695_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07951_ hold2516/X _07991_/A2 _07950_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _07951_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2906 _14633_/X vssd1 vssd1 vccd1 vccd1 _18109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2917 _17968_/Q vssd1 vssd1 vccd1 vccd1 hold2917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2928 _16204_/Q vssd1 vssd1 vccd1 vccd1 hold2928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2939 _14705_/X vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07882_ hold2254/X _07865_/B _07881_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _07882_/X
+ sky130_fd_sc_hd__o211a_1
X_09621_ _09933_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09552_ _09954_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09552_/X sky130_fd_sc_hd__or2_1
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ _08504_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _09483_/A hold634/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and3_1
XFILLER_0_19_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ hold2572/X _08433_/B _08433_/Y _08391_/A vssd1 vssd1 vccd1 vccd1 _08434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _12753_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _15814_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ hold2495/X _08336_/A2 _08295_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5510 _16768_/Q vssd1 vssd1 vccd1 vccd1 hold5510/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5521 _11026_/X vssd1 vssd1 vccd1 vccd1 _16832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5532 _16357_/Q vssd1 vssd1 vccd1 vccd1 hold5532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5543 _09808_/X vssd1 vssd1 vccd1 vccd1 _16426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5554 _16859_/Q vssd1 vssd1 vccd1 vccd1 hold5554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5565 _12052_/X vssd1 vssd1 vccd1 vccd1 _17174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4820 _17208_/Q vssd1 vssd1 vccd1 vccd1 hold4820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4831 _16788_/Q vssd1 vssd1 vccd1 vccd1 hold4831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5576 _16844_/Q vssd1 vssd1 vccd1 vccd1 hold5576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4842 hold5819/X vssd1 vssd1 vccd1 vccd1 hold4842/X sky130_fd_sc_hd__clkbuf_4
Xhold5587 _10678_/X vssd1 vssd1 vccd1 vccd1 _16716_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_86_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17343_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4853 _11716_/X vssd1 vssd1 vccd1 vccd1 _17062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5598 _16362_/Q vssd1 vssd1 vccd1 vccd1 hold5598/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4864 _16689_/Q vssd1 vssd1 vccd1 vccd1 hold4864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4875 _16932_/Q vssd1 vssd1 vccd1 vccd1 hold4875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4886 _09943_/X vssd1 vssd1 vccd1 vccd1 _16471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout320 _10515_/A vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__buf_2
Xhold4897 _17593_/Q vssd1 vssd1 vccd1 vccd1 hold4897/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17484_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout331 _10527_/A vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__buf_4
Xfanout342 _09369_/X vssd1 vssd1 vccd1 vccd1 _15483_/B sky130_fd_sc_hd__buf_4
Xfanout353 _08730_/X vssd1 vssd1 vccd1 vccd1 _08793_/S sky130_fd_sc_hd__buf_8
Xfanout364 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15221_/B sky130_fd_sc_hd__clkbuf_8
Xfanout375 _14966_/Y vssd1 vssd1 vccd1 vccd1 _15006_/B sky130_fd_sc_hd__buf_6
Xfanout386 _14784_/B vssd1 vssd1 vccd1 vccd1 _14786_/B sky130_fd_sc_hd__clkbuf_8
X_09819_ _09918_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__or2_1
Xfanout397 _14501_/Y vssd1 vssd1 vccd1 vccd1 _14554_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12830_ hold3044/X _12829_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__mux2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ hold3122/X _12760_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__mux2_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ hold895/X _14487_/B _14499_/X _14362_/A vssd1 vssd1 vccd1 vccd1 hold896/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12018_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__or2_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15489_/A _15480_/B _15480_/C _15480_/D vssd1 vssd1 vccd1 vccd1 _15480_/X
+ sky130_fd_sc_hd__or4_1
X_12692_ hold3050/X _12691_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__mux2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11652_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/X sky130_fd_sc_hd__or2_1
X_14431_ _15219_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__nand2_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ _17584_/CLK _17150_/D vssd1 vssd1 vccd1 vccd1 _17150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ _11670_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__or2_1
X_14362_ _14362_/A _14362_/B vssd1 vssd1 vccd1 vccd1 _17980_/D sky130_fd_sc_hd__and2_1
Xinput17 hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__clkbuf_2
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
X_16101_ _17525_/CLK _16101_/D vssd1 vssd1 vccd1 vccd1 hold620/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _10619_/A _10619_/B _10524_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _10525_/X
+ sky130_fd_sc_hd__o211a_1
X_13313_ hold1788/X hold4989/X _13793_/S vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__mux2_1
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
X_17081_ _17769_/CLK _17081_/D vssd1 vssd1 vccd1 vccd1 _17081_/Q sky130_fd_sc_hd__dfxtp_1
X_14293_ hold2664/X _14333_/A2 _14292_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14293_/X
+ sky130_fd_sc_hd__o211a_1
X_16032_ _17522_/CLK _16032_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
X_13244_ hold5309/X _13243_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ hold4127/X _10589_/B _10455_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10456_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _13183_/A1 _13173_/X _13174_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10387_ hold4565/X _10073_/B _10386_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12126_ _12267_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__or2_1
X_17983_ _18461_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
X_12057_ _12153_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__or2_1
X_16934_ _17877_/CLK _16934_/D vssd1 vssd1 vccd1 vccd1 _16934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ hold5536/X _11213_/B _11007_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__o211a_1
X_16865_ _18070_/CLK _16865_/D vssd1 vssd1 vccd1 vccd1 _16865_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _17697_/CLK _15816_/D vssd1 vssd1 vccd1 vccd1 _15816_/Q sky130_fd_sc_hd__dfxtp_1
X_16796_ _18060_/CLK _16796_/D vssd1 vssd1 vccd1 vccd1 _16796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _17686_/CLK _15747_/D vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ hold3104/X _12958_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_158_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15678_ _17170_/CLK _15678_/D vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17417_ _17419_/CLK _17417_/D vssd1 vssd1 vccd1 vccd1 _17417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14629_ hold2882/X _14666_/B _14628_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14629_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18397_ _18397_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _14728_/A hold2243/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__mux2_1
X_17348_ _17513_/CLK _17348_/D vssd1 vssd1 vccd1 vccd1 _17348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08081_ hold1257/X _08082_/B _08080_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17279_ _17279_/CLK _17279_/D vssd1 vssd1 vccd1 vccd1 _17279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4105 _16681_/Q vssd1 vssd1 vccd1 vccd1 hold4105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4116 _10999_/X vssd1 vssd1 vccd1 vccd1 _16823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4127 _16674_/Q vssd1 vssd1 vccd1 vccd1 hold4127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4138 _11365_/X vssd1 vssd1 vccd1 vccd1 _16945_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3404 _17134_/Q vssd1 vssd1 vccd1 vccd1 hold3404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4149 _16708_/Q vssd1 vssd1 vccd1 vccd1 hold4149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3415 _17349_/Q vssd1 vssd1 vccd1 vccd1 hold3415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3426 _17505_/Q vssd1 vssd1 vccd1 vccd1 hold3426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3437 _12527_/X vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08983_ hold251/X hold354/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__mux2_1
Xhold3448 _17436_/Q vssd1 vssd1 vccd1 vccd1 hold3448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2703 _18236_/Q vssd1 vssd1 vccd1 vccd1 hold2703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2714 _14522_/X vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3459 hold5856/X vssd1 vssd1 vccd1 vccd1 hold5857/A sky130_fd_sc_hd__buf_4
Xhold2725 _15773_/Q vssd1 vssd1 vccd1 vccd1 hold2725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2736 _18219_/Q vssd1 vssd1 vccd1 vccd1 hold2736/X sky130_fd_sc_hd__dlygate4sd3_1
X_07934_ _15557_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__or2_1
Xhold2747 _14759_/X vssd1 vssd1 vccd1 vccd1 _18170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _17909_/Q vssd1 vssd1 vccd1 vccd1 hold2758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 _17787_/Q vssd1 vssd1 vccd1 vccd1 hold2769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07865_ _15217_/A _07865_/B vssd1 vssd1 vccd1 vccd1 _07865_/Y sky130_fd_sc_hd__nand2_1
X_09604_ hold5524/X _10780_/A2 _09603_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _09604_/X
+ sky130_fd_sc_hd__o211a_1
X_07796_ _11155_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _07796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ hold5327/X _10028_/B _09534_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09535_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18378_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _09472_/C _09472_/D _09481_/B vssd1 vssd1 vccd1 vccd1 _09466_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ _15531_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__or2_1
X_09397_ hold5857/A _09342_/B _09342_/Y _09396_/X _12442_/A vssd1 vssd1 vccd1 vccd1
+ _09397_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _14511_/A hold977/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08279_ hold2568/X _08268_/B _08278_/X _12753_/A vssd1 vssd1 vccd1 vccd1 _08279_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6030 _16516_/Q vssd1 vssd1 vccd1 vccd1 hold6030/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6041 _18407_/Q vssd1 vssd1 vccd1 vccd1 hold6041/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10310_ hold2268/X hold3965/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__mux2_1
X_11290_ hold5739/X _11789_/B _11289_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5340 _16759_/Q vssd1 vssd1 vccd1 vccd1 hold5340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5351 _09745_/X vssd1 vssd1 vccd1 vccd1 _16405_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10241_ hold1905/X hold3976/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5362 _11593_/X vssd1 vssd1 vccd1 vccd1 _17021_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5373 _17011_/Q vssd1 vssd1 vccd1 vccd1 hold5373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5384 _09925_/X vssd1 vssd1 vccd1 vccd1 _16465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5395 _17081_/Q vssd1 vssd1 vccd1 vccd1 hold5395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4650 _11509_/X vssd1 vssd1 vccd1 vccd1 _16993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4661 _17251_/Q vssd1 vssd1 vccd1 vccd1 hold4661/X sky130_fd_sc_hd__dlygate4sd3_1
X_10172_ hold2218/X _16548_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__mux2_1
Xhold4672 _12076_/X vssd1 vssd1 vccd1 vccd1 _17182_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4683 _13729_/X vssd1 vssd1 vccd1 vccd1 _17696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4694 _17056_/Q vssd1 vssd1 vccd1 vccd1 hold4694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3960 _15490_/X vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14980_ _14980_/A _15012_/B vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__or2_1
Xhold3971 _13882_/Y vssd1 vssd1 vccd1 vccd1 _17747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3982 _10075_/Y vssd1 vssd1 vccd1 vccd1 _16515_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout150 _12836_/S vssd1 vssd1 vccd1 vccd1 _12848_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout161 _09494_/X vssd1 vssd1 vccd1 vccd1 _13808_/B sky130_fd_sc_hd__clkbuf_4
Xhold3993 _16887_/Q vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout172 _11617_/A2 vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__buf_4
X_13931_ _13931_/A hold403/X vssd1 vssd1 vccd1 vccd1 _17773_/D sky130_fd_sc_hd__and2_1
Xfanout183 _09494_/X vssd1 vssd1 vccd1 vccd1 _10852_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout194 _12374_/B vssd1 vssd1 vccd1 vccd1 _13844_/B sky130_fd_sc_hd__buf_4
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16650_ _18353_/CLK _16650_/D vssd1 vssd1 vccd1 vccd1 _16650_/Q sky130_fd_sc_hd__dfxtp_1
X_13862_ _17741_/Q _13862_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _17217_/CLK _15601_/D vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfxtp_1
X_12813_ _12813_/A _12813_/B vssd1 vssd1 vccd1 vccd1 _17447_/D sky130_fd_sc_hd__and2_1
X_16581_ _18235_/CLK _16581_/D vssd1 vssd1 vccd1 vccd1 _16581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13793_ hold2639/X hold3324/X _13793_/S vssd1 vssd1 vccd1 vccd1 _13794_/B sky130_fd_sc_hd__mux2_1
X_18320_ _18390_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ hold1346/X _15547_/B _15531_/X _12825_/A vssd1 vssd1 vccd1 vccd1 _15532_/X
+ sky130_fd_sc_hd__o211a_1
X_12744_ _12753_/A _12744_/B vssd1 vssd1 vccd1 vccd1 _17424_/D sky130_fd_sc_hd__and2_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18373_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15481_/A1 _15455_/X _15462_/X _15481_/B1 _18422_/Q vssd1 vssd1 vccd1 vccd1
+ _15463_/X sky130_fd_sc_hd__a32o_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12675_ _12876_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _17401_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17202_ _17266_/CLK _17202_/D vssd1 vssd1 vccd1 vccd1 _17202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ hold2491/X hold209/X _14413_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14414_/X
+ sky130_fd_sc_hd__o211a_1
X_18182_ _18206_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
X_11626_ hold4631/X _12299_/B _11625_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11626_/X
+ sky130_fd_sc_hd__o211a_1
X_15394_ _15394_/A _15394_/B vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17133_ _17252_/CLK _17133_/D vssd1 vssd1 vccd1 vccd1 _17133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14345_ _14740_/A hold2596/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14346_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ hold4101/X _11747_/B _11556_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ hold1531/X _16660_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10509_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _17257_/CLK _17064_/D vssd1 vssd1 vccd1 vccd1 _17064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold609 hold609/A vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__buf_6
X_11488_ hold5540/X _12338_/B _11487_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11488_/X
+ sky130_fd_sc_hd__o211a_1
X_14276_ _14330_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ _18422_/CLK _16015_/D vssd1 vssd1 vccd1 vccd1 _16015_/Q sky130_fd_sc_hd__dfxtp_1
X_10439_ hold2180/X _16637_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ _13226_/X hold5236/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13227_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13158_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__or2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ hold4655/X _12299_/B _12108_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _12109_/X
+ sky130_fd_sc_hd__o211a_1
X_13089_ _13089_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__and2_1
X_17966_ _18054_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1309 _17866_/Q vssd1 vssd1 vccd1 vccd1 hold1309/X sky130_fd_sc_hd__dlygate4sd3_1
X_16917_ _17829_/CLK _16917_/D vssd1 vssd1 vccd1 vccd1 _16917_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _17897_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16848_ _18052_/CLK _16848_/D vssd1 vssd1 vccd1 vccd1 _16848_/Q sky130_fd_sc_hd__dfxtp_1
X_16779_ _18305_/CLK _16779_/D vssd1 vssd1 vccd1 vccd1 _16779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09320_ hold2123/X _09325_/B _09319_/Y _15504_/A vssd1 vssd1 vccd1 vccd1 _09320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ _15527_/A hold2455/X _09283_/S vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18449_ _18450_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
X_08202_ hold1765/X _08213_/B _08201_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _08202_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ hold892/X _09230_/B vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _15705_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ hold949/X _08094_/B vssd1 vssd1 vccd1 vccd1 _08064_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3201 _17478_/Q vssd1 vssd1 vccd1 vccd1 hold3201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3212 _17656_/Q vssd1 vssd1 vccd1 vccd1 hold3212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3223 _16880_/Q vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3234 _16663_/Q vssd1 vssd1 vccd1 vccd1 hold3234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2500 _14675_/X vssd1 vssd1 vccd1 vccd1 _18130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3245 _12557_/X vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3256 _13705_/X vssd1 vssd1 vccd1 vccd1 _17688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2511 _16171_/Q vssd1 vssd1 vccd1 vccd1 hold2511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3267 _17132_/Q vssd1 vssd1 vccd1 vccd1 hold3267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 _15644_/Q vssd1 vssd1 vccd1 vccd1 hold2522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 _15013_/X vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08966_ _09063_/A hold258/X vssd1 vssd1 vccd1 vccd1 _16100_/D sky130_fd_sc_hd__and2_1
Xhold3278 _13768_/X vssd1 vssd1 vccd1 vccd1 _17709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3289 _17465_/Q vssd1 vssd1 vccd1 vccd1 hold3289/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2544 _16169_/Q vssd1 vssd1 vccd1 vccd1 hold2544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1810 _14599_/X vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 _15877_/Q vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 _08324_/X vssd1 vssd1 vccd1 vccd1 _15795_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07917_ hold1359/X _07918_/B _07916_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07917_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2566 _16260_/Q vssd1 vssd1 vccd1 vccd1 hold2566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2577 _15076_/X vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1832 _15605_/Q vssd1 vssd1 vccd1 vccd1 hold1832/X sky130_fd_sc_hd__dlygate4sd3_1
X_08897_ _12402_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _16066_/D sky130_fd_sc_hd__and2_1
Xhold2588 _15762_/Q vssd1 vssd1 vccd1 vccd1 hold2588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 _15812_/Q vssd1 vssd1 vccd1 vccd1 hold1843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1854 _18453_/Q vssd1 vssd1 vccd1 vccd1 hold1854/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_314_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold2599 _16188_/Q vssd1 vssd1 vccd1 vccd1 hold2599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1865 _08416_/X vssd1 vssd1 vccd1 vccd1 _15838_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1876 _15711_/Q vssd1 vssd1 vccd1 vccd1 hold1876/X sky130_fd_sc_hd__dlygate4sd3_1
X_07848_ hold2072/X _07869_/B _07847_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _07848_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1887 _18089_/Q vssd1 vssd1 vccd1 vccd1 hold1887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1898 _16238_/Q vssd1 vssd1 vccd1 vccd1 hold1898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ hold1899/X _13110_/A _09998_/C vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ hold1665/X _16754_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__mux2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09456_/D _09449_/B vssd1 vssd1 vccd1 vccd1 _16309_/D sky130_fd_sc_hd__nor2_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ _17323_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ hold2723/X _16961_/Q _12341_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__mux2_1
X_12391_ hold41/X hold309/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14130_ hold747/X _14138_/B vssd1 vssd1 vccd1 vccd1 hold748/A sky130_fd_sc_hd__or2_1
X_11342_ hold904/X _16938_/Q _11726_/C vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17852_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14061_ hold2975/X _14105_/A2 _14060_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _14061_/X
+ sky130_fd_sc_hd__o211a_1
X_11273_ hold1239/X hold5233/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5170 hold6030/X vssd1 vssd1 vccd1 vccd1 hold5170/X sky130_fd_sc_hd__clkbuf_2
X_10224_ _10554_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__or2_1
Xhold5181 hold5833/X vssd1 vssd1 vccd1 vccd1 hold5181/X sky130_fd_sc_hd__buf_4
X_13012_ hold683/X _13003_/Y _13011_/X _12936_/A vssd1 vssd1 vccd1 vccd1 hold684/A
+ sky130_fd_sc_hd__o211a_1
Xhold5192 _15463_/X vssd1 vssd1 vccd1 vccd1 _15464_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4480 _17604_/Q vssd1 vssd1 vccd1 vccd1 hold4480/X sky130_fd_sc_hd__dlygate4sd3_1
X_17820_ _17852_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4491 _12175_/X vssd1 vssd1 vccd1 vccd1 _17215_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10155_ _10521_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__or2_1
XFILLER_0_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3790 _16912_/Q vssd1 vssd1 vccd1 vccd1 hold3790/X sky130_fd_sc_hd__dlygate4sd3_1
X_17751_ _17751_/CLK _17751_/D vssd1 vssd1 vccd1 vccd1 _17751_/Q sky130_fd_sc_hd__dfxtp_1
X_14963_ hold1373/X _14946_/B _14962_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14963_/X
+ sky130_fd_sc_hd__o211a_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _10563_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16702_ _18228_/CLK _16702_/D vssd1 vssd1 vccd1 vccd1 _16702_/Q sky130_fd_sc_hd__dfxtp_1
X_13914_ hold747/X _17765_/Q hold244/X vssd1 vssd1 vccd1 vccd1 hold753/A sky130_fd_sc_hd__mux2_1
X_17682_ _17747_/CLK _17682_/D vssd1 vssd1 vccd1 vccd1 _17682_/Q sky130_fd_sc_hd__dfxtp_1
X_14894_ _15233_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14894_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16633_ _18095_/CLK _16633_/D vssd1 vssd1 vccd1 vccd1 _16633_/Q sky130_fd_sc_hd__dfxtp_1
X_13845_ hold3902/X _13749_/A _13844_/X vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16564_ _18218_/CLK _16564_/D vssd1 vssd1 vccd1 vccd1 _16564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13776_/X sky130_fd_sc_hd__or2_1
X_10988_ hold1399/X _16820_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _10989_/B sky130_fd_sc_hd__mux2_1
X_18303_ _18337_/CLK hold951/X vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15515_ _15515_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15515_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12727_ hold2378/X hold3468/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16495_ _18416_/CLK _16495_/D vssd1 vssd1 vccd1 vccd1 _16495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18234_ _18236_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
X_15446_ _17320_/Q _09357_/A _15446_/B1 hold277/X vssd1 vssd1 vccd1 vccd1 _15446_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ hold1480/X _17397_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18165_ _18183_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
X_11609_ hold2172/X _17027_/Q _12341_/C vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__mux2_1
X_15377_ hold642/X _15479_/A2 _09386_/D hold533/X _15376_/X vssd1 vssd1 vccd1 vccd1
+ _15382_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_26_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ hold2165/X _17374_/Q _12589_/S vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _17742_/CLK _17116_/D vssd1 vssd1 vccd1 vccd1 _17116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _15169_/A _14334_/B vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__or2_1
X_18096_ _18218_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold406 input27/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold417 hold417/A vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 hold570/X vssd1 vssd1 vccd1 vccd1 hold571/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _17895_/CLK _17047_/D vssd1 vssd1 vccd1 vccd1 _17047_/Q sky130_fd_sc_hd__dfxtp_1
X_14259_ hold2742/X _14272_/B _14258_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14259_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 hold1030/X vssd1 vssd1 vccd1 vccd1 hold1031/A sky130_fd_sc_hd__buf_6
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 hold573/X vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__buf_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ hold126/X hold446/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _08018_/X vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _14179_/X vssd1 vssd1 vccd1 vccd1 _17892_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ hold53/X hold579/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__mux2_1
Xhold1128 _15861_/Q vssd1 vssd1 vccd1 vccd1 hold1128/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _18047_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1139 _14167_/X vssd1 vssd1 vccd1 vccd1 _17886_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08682_ _08970_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _15962_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ _14984_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09234_ _12849_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _16228_/D sky130_fd_sc_hd__and2_1
XFILLER_0_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09165_ hold1840/X _09177_/A2 _09164_/Y _12909_/A vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__o211a_1
X_08116_ _14246_/A hold2766/X hold196/X vssd1 vssd1 vccd1 vccd1 _08117_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ _15103_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08047_ hold624/A hold279/X hold606/A hold298/X vssd1 vssd1 vccd1 vccd1 _14627_/A
+ sky130_fd_sc_hd__or4bb_4
Xhold940 hold940/A vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold951 hold951/A vssd1 vssd1 vccd1 vccd1 hold951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3020 _17383_/Q vssd1 vssd1 vccd1 vccd1 hold3020/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3031 _17389_/Q vssd1 vssd1 vccd1 vccd1 hold3031/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3042 _17488_/Q vssd1 vssd1 vccd1 vccd1 hold3042/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3053 _12788_/X vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3064 _12845_/X vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__dlygate4sd3_1
X_09998_ _16490_/Q _09998_/B _09998_/C vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__and3_1
Xhold3075 _12623_/X vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2330 _17847_/Q vssd1 vssd1 vccd1 vccd1 hold2330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2341 _12836_/X vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3086 _17386_/Q vssd1 vssd1 vccd1 vccd1 hold3086/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2352 _15772_/Q vssd1 vssd1 vccd1 vccd1 hold2352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3097 _17502_/Q vssd1 vssd1 vccd1 vccd1 hold3097/X sky130_fd_sc_hd__dlygate4sd3_1
X_08949_ hold47/X hold552/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__mux2_1
Xhold2363 _18147_/Q vssd1 vssd1 vccd1 vccd1 hold2363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2374 _16167_/Q vssd1 vssd1 vccd1 vccd1 hold2374/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _15831_/Q vssd1 vssd1 vccd1 vccd1 hold1640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 _09225_/X vssd1 vssd1 vccd1 vccd1 _16224_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1651 _08257_/X vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2396 _15717_/Q vssd1 vssd1 vccd1 vccd1 hold2396/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ hold2469/X hold3362/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__mux2_1
Xhold1662 _14171_/X vssd1 vssd1 vccd1 vccd1 _17888_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1673 _18140_/Q vssd1 vssd1 vccd1 vccd1 hold1673/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1684 _18329_/Q vssd1 vssd1 vccd1 vccd1 hold1684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1695 _07893_/X vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10911_ _11103_/A _10911_/B vssd1 vssd1 vccd1 vccd1 _10911_/X sky130_fd_sc_hd__or2_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ hold1848/X hold3828/X _12377_/C vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__mux2_1
X_13630_ hold4167/X _13829_/B _13629_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13630_/X
+ sky130_fd_sc_hd__o211a_1
X_10842_ _11031_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ hold5132/X _13847_/B _13560_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10773_ _11136_/A _10773_/B vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__or2_1
X_15300_ hold522/X _15486_/A2 _15446_/B1 hold576/X vssd1 vssd1 vccd1 vccd1 _15300_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ _09342_/A hold2175/X _07802_/Y _12511_/X vssd1 vssd1 vccd1 vccd1 _12512_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16280_ _17751_/CLK _16280_/D vssd1 vssd1 vccd1 vccd1 _16280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13492_ hold5146/X _13883_/B _13491_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15231_ _15231_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ hold291/X hold338/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ hold1267/X _15161_/B _15161_/Y _15070_/A vssd1 vssd1 vccd1 vccd1 _15162_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12374_ _12374_/A _12374_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__and3_1
X_14113_ hold983/X hold587/X _14112_/X _13913_/A vssd1 vssd1 vccd1 vccd1 hold984/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11325_ _11649_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__or2_1
X_15093_ hold883/X _15123_/B vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044_ _14330_/A _14050_/B vssd1 vssd1 vccd1 vccd1 _14044_/X sky130_fd_sc_hd__or2_1
X_11256_ _11640_/A _11256_/B vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_236_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17745_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ hold4188/X _10631_/B _10206_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10207_/X
+ sky130_fd_sc_hd__o211a_1
X_11187_ hold3784/X _11097_/A _11186_/X vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17803_ _17855_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_1
X_10138_ hold4295/X _10643_/B _10137_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15995_ _18409_/CLK _15995_/D vssd1 vssd1 vccd1 vccd1 hold452/A sky130_fd_sc_hd__dfxtp_1
X_17734_ _17734_/CLK _17734_/D vssd1 vssd1 vccd1 vccd1 _17734_/Q sky130_fd_sc_hd__dfxtp_1
X_10069_ _10588_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10069_/Y sky130_fd_sc_hd__nor2_1
X_14946_ _15215_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _17697_/CLK _17665_/D vssd1 vssd1 vccd1 vccd1 _17665_/Q sky130_fd_sc_hd__dfxtp_1
X_14877_ hold989/X _14880_/B _14876_/Y _14877_/C1 vssd1 vssd1 vccd1 vccd1 hold990/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16616_ _18265_/CLK _16616_/D vssd1 vssd1 vccd1 vccd1 _16616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13828_ _13864_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13828_/Y sky130_fd_sc_hd__nor2_1
X_17596_ _17724_/CLK _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16547_ _18233_/CLK _16547_/D vssd1 vssd1 vccd1 vccd1 _16547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13759_ hold4943/X _13859_/B _13758_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16478_ _18391_/CLK _16478_/D vssd1 vssd1 vccd1 vccd1 _16478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18217_ _18217_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15429_ hold416/X _09386_/A _15427_/X vssd1 vssd1 vccd1 vccd1 _15432_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18148_ _18265_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5906 _17530_/Q vssd1 vssd1 vccd1 vccd1 hold5906/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5917 _17540_/Q vssd1 vssd1 vccd1 vccd1 hold5917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5928 _17542_/Q vssd1 vssd1 vccd1 vccd1 hold5928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 input30/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 hold20/X vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__buf_4
Xhold5939 hold5996/X vssd1 vssd1 vccd1 vccd1 hold5939/X sky130_fd_sc_hd__buf_1
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _18319_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold812/X vssd1 vssd1 vccd1 vccd1 hold813/A sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _09987_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout705 _08887_/A vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__buf_2
XFILLER_0_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout716 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__buf_4
X_09852_ _09948_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__or2_1
Xfanout727 _08585_/A vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 fanout842/X vssd1 vssd1 vccd1 vccd1 _08585_/A sky130_fd_sc_hd__clkbuf_8
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _12142_/C1 vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__buf_4
X_08803_ _08868_/B _12380_/B _13046_/D vssd1 vssd1 vccd1 vccd1 _08866_/S sky130_fd_sc_hd__or3_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09975_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _15482_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _15987_/D sky130_fd_sc_hd__and2_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _14980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ hold23/X hold325/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08666_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _13043_/C _17518_/Q vssd1 vssd1 vccd1 vccd1 _13034_/D sky130_fd_sc_hd__and2_2
XFILLER_0_152_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09217_ hold2018/X _09216_/B _09216_/Y _15534_/C1 vssd1 vssd1 vccd1 vccd1 _09217_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ _15531_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ hold2451/X _09119_/A2 _09078_/X _12996_/A vssd1 vssd1 vccd1 vccd1 _09079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _11204_/A _11210_/B _11109_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11110_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _12282_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__or2_1
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__buf_12
Xhold781 hold781/A vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold792 input4/X vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ hold5623/X _11156_/B _11040_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _11041_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _15104_/X vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2171 _14193_/X vssd1 vssd1 vccd1 vccd1 _17899_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _15193_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__or2_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 _15811_/Q vssd1 vssd1 vccd1 vccd1 hold2182/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _17647_/CLK _15780_/D vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2193 _17803_/Q vssd1 vssd1 vccd1 vccd1 hold2193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ hold3424/X _12991_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__mux2_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1470 _14767_/X vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ hold2293/X _14718_/B _14730_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _14731_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1481 _15540_/X vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _12243_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__or2_1
Xhold1492 _14135_/X vssd1 vssd1 vccd1 vccd1 _17871_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17456_/CLK _17450_/D vssd1 vssd1 vccd1 vccd1 _17450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _15217_/A _14666_/B vssd1 vssd1 vccd1 vccd1 _14662_/Y sky130_fd_sc_hd__nand2_1
X_11874_ _12267_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__or2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _18378_/CLK _16401_/D vssd1 vssd1 vccd1 vccd1 _16401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ hold1041/X hold3251/X _13805_/C vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17381_ _17464_/CLK _17381_/D vssd1 vssd1 vccd1 vccd1 _17381_/Q sky130_fd_sc_hd__dfxtp_1
X_10825_ hold5733/X _11222_/B _10824_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10825_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ hold2683/X _14612_/B _14592_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16332_ _18424_/CLK _16332_/D vssd1 vssd1 vccd1 vccd1 _16332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13544_ _15820_/Q _17635_/Q _13832_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10756_ hold4341/X _11732_/B _10755_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _10756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16263_ _17494_/CLK _16263_/D vssd1 vssd1 vccd1 vccd1 _16263_/Q sky130_fd_sc_hd__dfxtp_1
X_13475_ hold1328/X hold5168/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__mux2_1
X_10687_ hold4131/X _11201_/B _10686_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _10687_/X
+ sky130_fd_sc_hd__o211a_1
X_18002_ _18034_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ hold1317/X _15221_/B _15213_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _15214_/X
+ sky130_fd_sc_hd__o211a_1
X_12426_ _12426_/A hold711/X vssd1 vssd1 vccd1 vccd1 _17306_/D sky130_fd_sc_hd__and2_1
XFILLER_0_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _17480_/CLK _16194_/D vssd1 vssd1 vccd1 vccd1 _16194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15145_ _15199_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12357_ hold3897/X _12267_/A _12356_/X vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11308_ hold5494/X _11783_/B _11307_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 _11308_/X
+ sky130_fd_sc_hd__o211a_1
X_15076_ hold2576/X _15113_/B _15075_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _15076_/X
+ sky130_fd_sc_hd__o211a_1
X_12288_ _13797_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__or2_1
X_14027_ hold2616/X _14040_/B _14026_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14027_/X
+ sky130_fd_sc_hd__o211a_1
X_11239_ hold3382/X _12299_/B _11238_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _11239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _18425_/CLK _15978_/D vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ hold1571/X _14952_/B _14928_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _14929_/X
+ sky130_fd_sc_hd__o211a_1
X_17717_ _17749_/CLK _17717_/D vssd1 vssd1 vccd1 vccd1 _17717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ _14218_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08450_/X sky130_fd_sc_hd__or2_1
X_17648_ _17739_/CLK _17648_/D vssd1 vssd1 vccd1 vccd1 _17648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _15822_/D sky130_fd_sc_hd__and2_1
X_17579_ _17734_/CLK _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09002_ hold68/X hold646/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5703 _16878_/Q vssd1 vssd1 vccd1 vccd1 hold5703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5714 _11695_/X vssd1 vssd1 vccd1 vccd1 _17055_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_158_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5725 _16770_/Q vssd1 vssd1 vccd1 vccd1 hold5725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5736 _11377_/X vssd1 vssd1 vccd1 vccd1 _16949_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5747 _16950_/Q vssd1 vssd1 vccd1 vccd1 hold5747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5758 output97/X vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_12
Xhold5769 hold5913/X vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__buf_1
Xfanout502 _10568_/C vssd1 vssd1 vccd1 vccd1 _10565_/C sky130_fd_sc_hd__clkbuf_8
X_09904_ hold5552/X _09998_/B _09903_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09904_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout513 fanout523/X vssd1 vssd1 vccd1 vccd1 _10067_/C sky130_fd_sc_hd__buf_4
Xfanout524 _09340_/X vssd1 vssd1 vccd1 vccd1 _15490_/B1 sky130_fd_sc_hd__buf_6
Xfanout535 _09177_/A2 vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__buf_4
Xfanout546 _08448_/Y vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__clkbuf_8
X_09835_ hold4059/X _10001_/B _09834_/X _15208_/C1 vssd1 vssd1 vccd1 vccd1 _09835_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout557 _08228_/Y vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__clkbuf_8
Xfanout568 _07993_/Y vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__clkbuf_8
Xfanout579 _14610_/B vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__clkbuf_8
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ hold5492/X _10013_/B _09765_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09766_/X
+ sky130_fd_sc_hd__o211a_1
X_08717_ hold65/X hold132/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08718_/B sky130_fd_sc_hd__mux2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ hold5476/X _10016_/B _09696_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09697_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08648_ _13002_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _15946_/D sky130_fd_sc_hd__and2_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _12438_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _15913_/D sky130_fd_sc_hd__and2_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _16694_/Q _10610_/B _10610_/C vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11590_ hold4601/X _12323_/B _11589_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11590_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ hold2445/X hold3271/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13260_ hold5447/X _13259_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__mux2_2
X_10472_ hold1688/X _16648_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _12305_/A _12302_/B _12210_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _12211_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ _13311_/A1 _13189_/X _13190_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12142_ hold3444/X _12347_/B _12141_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _12142_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12073_ hold4990/X _13871_/B _12072_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _12073_/X
+ sky130_fd_sc_hd__o211a_1
X_16950_ _17798_/CLK _16950_/D vssd1 vssd1 vccd1 vccd1 _16950_/Q sky130_fd_sc_hd__dfxtp_1
X_15901_ _17345_/CLK _15901_/D vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__dfxtp_1
X_11024_ hold1748/X _16832_/Q _11216_/C vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__mux2_1
X_16881_ _18052_/CLK _16881_/D vssd1 vssd1 vccd1 vccd1 _16881_/Q sky130_fd_sc_hd__dfxtp_1
X_15832_ _17722_/CLK _15832_/D vssd1 vssd1 vccd1 vccd1 _15832_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _17747_/CLK _15763_/D vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _14364_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _17501_/D sky130_fd_sc_hd__and2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14714_ _15000_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14714_/Y sky130_fd_sc_hd__nand2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17502_ _17503_/CLK _17502_/D vssd1 vssd1 vccd1 vccd1 _17502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ hold3242/X _12302_/B _11925_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15694_ _17262_/CLK _15694_/D vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17435_/CLK _17433_/D vssd1 vssd1 vccd1 vccd1 _17433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ hold2139/X _14664_/B _14644_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _14645_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ hold4765/X _11798_/B _11856_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11857_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17364_ _17487_/CLK _17364_/D vssd1 vssd1 vccd1 vccd1 _17364_/Q sky130_fd_sc_hd__dfxtp_1
X_10808_ hold2564/X hold5596/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
X_14576_ hold756/X _14624_/B vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _12331_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11788_/Y sky130_fd_sc_hd__nor2_1
X_16315_ _17503_/CLK _16315_/D vssd1 vssd1 vccd1 vccd1 _16315_/Q sky130_fd_sc_hd__dfxtp_1
X_13527_ _13800_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__or2_1
X_17295_ _18411_/CLK _17295_/D vssd1 vssd1 vccd1 vccd1 hold561/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ hold1870/X hold3705/X _11219_/C vssd1 vssd1 vccd1 vccd1 _10740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16246_ _17666_/CLK hold337/X vssd1 vssd1 vccd1 vccd1 _16246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _13764_/A _13458_/B vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_251_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17647_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12409_ hold71/X hold353/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__mux2_1
X_16177_ _18441_/CLK hold974/X vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__dfxtp_1
X_13389_ _13758_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput105 _17524_/Q vssd1 vssd1 vccd1 vccd1 io_out sky130_fd_sc_hd__buf_12
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4309 _16477_/Q vssd1 vssd1 vccd1 vccd1 hold4309/X sky130_fd_sc_hd__dlygate4sd3_1
Xoutput116 hold5865/X vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_12
Xoutput127 hold5851/X vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_12
Xoutput138 hold5848/X vssd1 vssd1 vccd1 vccd1 hold5849/A sky130_fd_sc_hd__buf_6
X_15128_ hold607/X hold656/X vssd1 vssd1 vccd1 vccd1 _15149_/B sky130_fd_sc_hd__or2_4
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3608 _11148_/Y vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3619 _16536_/Q vssd1 vssd1 vccd1 vccd1 hold3619/X sky130_fd_sc_hd__buf_1
X_15059_ hold173/X hold362/X hold302/X vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__mux2_1
X_07950_ _14854_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07950_/X sky130_fd_sc_hd__or2_1
Xhold2907 _18142_/Q vssd1 vssd1 vccd1 vccd1 hold2907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 _14337_/X vssd1 vssd1 vccd1 vccd1 _17968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2929 _09185_/X vssd1 vssd1 vccd1 vccd1 _16204_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07881_ _15559_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07881_/X sky130_fd_sc_hd__or2_1
X_09620_ hold1595/X hold5338/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__mux2_1
X_09551_ hold822/X _13198_/A _10055_/C vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__mux2_1
X_08502_ hold624/A hold298/X hold606/A hold279/X vssd1 vssd1 vccd1 vccd1 _14897_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09482_ _09483_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09484_/C sky130_fd_sc_hd__or2_1
X_08433_ _14774_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ _15533_/A hold2093/X hold122/X vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ _14854_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08295_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5500 _16948_/Q vssd1 vssd1 vccd1 vccd1 hold5500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5511 _10738_/X vssd1 vssd1 vccd1 vccd1 _16736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5522 _17267_/Q vssd1 vssd1 vccd1 vccd1 hold5522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5533 _09505_/X vssd1 vssd1 vccd1 vccd1 _16325_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5544 _16489_/Q vssd1 vssd1 vccd1 vccd1 hold5544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4810 _12205_/X vssd1 vssd1 vccd1 vccd1 _17225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5555 _11011_/X vssd1 vssd1 vccd1 vccd1 _16827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5566 _16372_/Q vssd1 vssd1 vccd1 vccd1 hold5566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4821 _12058_/X vssd1 vssd1 vccd1 vccd1 _17176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4832 _16680_/Q vssd1 vssd1 vccd1 vccd1 hold4832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5577 _10966_/X vssd1 vssd1 vccd1 vccd1 _16812_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4843 _15273_/X vssd1 vssd1 vccd1 vccd1 _15274_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5588 _16478_/Q vssd1 vssd1 vccd1 vccd1 hold5588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4854 _16965_/Q vssd1 vssd1 vccd1 vccd1 hold4854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5599 _09520_/X vssd1 vssd1 vccd1 vccd1 _16330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4865 _17202_/Q vssd1 vssd1 vccd1 vccd1 hold4865/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4876 _11230_/X vssd1 vssd1 vccd1 vccd1 _16900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout310 _09948_/A vssd1 vssd1 vccd1 vccd1 _09924_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout321 _10515_/A vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__buf_4
Xhold4887 _17068_/Q vssd1 vssd1 vccd1 vccd1 hold4887/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout332 _10527_/A vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__buf_4
Xhold4898 _13324_/X vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout343 _09369_/X vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__clkbuf_4
Xfanout354 _08721_/S vssd1 vssd1 vccd1 vccd1 _08727_/S sky130_fd_sc_hd__buf_8
Xfanout365 _15181_/Y vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__clkbuf_8
Xfanout376 _14966_/Y vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__clkbuf_8
X_09818_ _18343_/Q _16430_/Q _09893_/S vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__mux2_1
Xfanout387 _14734_/Y vssd1 vssd1 vccd1 vccd1 _14774_/B sky130_fd_sc_hd__buf_8
Xfanout398 _14479_/B vssd1 vssd1 vccd1 vccd1 _14499_/B sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_55_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17494_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09749_ hold1277/X hold4528/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12760_ hold2678/X _17431_/Q _12814_/S vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ hold2758/X hold3351/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__mux2_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ hold2540/X _17408_/Q _12844_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ hold1925/X _14433_/B _14429_/Y _12984_/A vssd1 vssd1 vccd1 vccd1 _14430_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ hold1138/X _17038_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14988_/A hold2456/X hold275/X vssd1 vssd1 vccd1 vccd1 _14362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ hold1077/X _17015_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__mux2_1
Xinput18 input18/A vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
X_16100_ _17300_/CLK _16100_/D vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13312_ _13305_/X _13311_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__o21a_1
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or2_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17080_ _17903_/CLK _17080_/D vssd1 vssd1 vccd1 vccd1 _17080_/Q sky130_fd_sc_hd__dfxtp_1
X_14292_ _14972_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14292_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _17323_/CLK _16031_/D vssd1 vssd1 vccd1 vccd1 hold538/A sky130_fd_sc_hd__dfxtp_1
X_13243_ _13242_/X _16923_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__mux2_1
X_10455_ _10551_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13174_ _13174_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__or2_1
X_10386_ _10506_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ hold2392/X _17199_/Q _12356_/C vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__mux2_1
X_17982_ _18305_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
X_12056_ hold2145/X hold4639/X _12152_/S vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__mux2_1
X_16933_ _17877_/CLK _16933_/D vssd1 vssd1 vccd1 vccd1 _16933_/Q sky130_fd_sc_hd__dfxtp_1
X_11007_ _11103_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__or2_1
XFILLER_0_189_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16864_ _18067_/CLK _16864_/D vssd1 vssd1 vccd1 vccd1 _16864_/Q sky130_fd_sc_hd__dfxtp_1
X_15815_ _17726_/CLK _15815_/D vssd1 vssd1 vccd1 vccd1 _15815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16795_ _18054_/CLK _16795_/D vssd1 vssd1 vccd1 vccd1 _16795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15746_ _17749_/CLK _15746_/D vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ hold1482/X hold3084/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11909_ hold2646/X _17127_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15677_ _17900_/CLK _15677_/D vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfxtp_1
X_12889_ hold2332/X hold3018/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ _15129_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14628_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17416_ _17419_/CLK _17416_/D vssd1 vssd1 vccd1 vccd1 _17416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18396_ _18396_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17347_ _17531_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 _17347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14559_ _15129_/A _14557_/Y hold1802/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14559_/X
+ sky130_fd_sc_hd__o211a_1
X_08080_ _15539_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08080_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17278_ _17584_/CLK _17278_/D vssd1 vssd1 vccd1 vccd1 _17278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _17439_/CLK _16229_/D vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4106 _10477_/X vssd1 vssd1 vccd1 vccd1 _16649_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4117 _17655_/Q vssd1 vssd1 vccd1 vccd1 hold4117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4128 _10456_/X vssd1 vssd1 vccd1 vccd1 _16642_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4139 _17602_/Q vssd1 vssd1 vccd1 vccd1 hold4139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3405 _11836_/X vssd1 vssd1 vccd1 vccd1 _17102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3416 _17710_/Q vssd1 vssd1 vccd1 vccd1 hold3416/X sky130_fd_sc_hd__dlygate4sd3_1
X_08982_ _15284_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _16108_/D sky130_fd_sc_hd__and2_1
Xhold3427 _17138_/Q vssd1 vssd1 vccd1 vccd1 hold3427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3438 _17354_/Q vssd1 vssd1 vccd1 vccd1 hold3438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3449 _12779_/X vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2704 _14895_/X vssd1 vssd1 vccd1 vccd1 _18236_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2715 _17952_/Q vssd1 vssd1 vccd1 vccd1 hold2715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2726 _08277_/X vssd1 vssd1 vccd1 vccd1 _15773_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07933_ hold2113/X _07924_/B _07932_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _07933_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2737 _14861_/X vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2748 _18385_/Q vssd1 vssd1 vccd1 vccd1 hold2748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 _14213_/X vssd1 vssd1 vccd1 vccd1 _17909_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07864_ hold2102/X _07869_/B _07863_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 _07864_/X
+ sky130_fd_sc_hd__o211a_1
X_09603_ _11067_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07795_ _18461_/Q hold1119/X _09342_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _07795_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09534_ _09918_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09472_/D _09465_/B vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_176_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08416_ hold1864/X _08440_/A2 _08415_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08416_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _09386_/B _09369_/B _18460_/Q vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_173_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18158_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08347_ _08391_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__and2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_102_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _16128_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08278_ _15557_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__or2_1
Xhold6020 data_in[6] vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6031 la_data_in[4] vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5330 _10747_/X vssd1 vssd1 vccd1 vccd1 _16739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10240_ hold4242/X _10640_/B _10239_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10240_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5341 _10711_/X vssd1 vssd1 vccd1 vccd1 _16727_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5352 _16453_/Q vssd1 vssd1 vccd1 vccd1 hold5352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5363 _16366_/Q vssd1 vssd1 vccd1 vccd1 hold5363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5374 _11467_/X vssd1 vssd1 vccd1 vccd1 _16979_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5385 _16468_/Q vssd1 vssd1 vccd1 vccd1 hold5385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4640 _11962_/X vssd1 vssd1 vccd1 vccd1 _17144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10171_ hold3206/X _10649_/B _10170_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _10171_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4651 _17636_/Q vssd1 vssd1 vccd1 vccd1 hold4651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5396 _11677_/X vssd1 vssd1 vccd1 vccd1 _17049_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4662 _12187_/X vssd1 vssd1 vccd1 vccd1 _17219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4673 _17680_/Q vssd1 vssd1 vccd1 vccd1 hold4673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4684 _17228_/Q vssd1 vssd1 vccd1 vccd1 hold4684/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3950 _17099_/Q vssd1 vssd1 vccd1 vccd1 hold3950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4695 _11602_/X vssd1 vssd1 vccd1 vccd1 _17024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3961 _16874_/Q vssd1 vssd1 vccd1 vccd1 hold3961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout151 _12836_/S vssd1 vssd1 vccd1 vccd1 _12677_/S sky130_fd_sc_hd__clkbuf_8
Xhold3972 _16658_/Q vssd1 vssd1 vccd1 vccd1 hold3972/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout162 _12302_/B vssd1 vssd1 vccd1 vccd1 _13811_/B sky130_fd_sc_hd__buf_4
Xhold3983 _16782_/Q vssd1 vssd1 vccd1 vccd1 hold3983/X sky130_fd_sc_hd__dlygate4sd3_1
X_13930_ hold335/X hold402/X hold244/X vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__mux2_1
Xhold3994 _11095_/X vssd1 vssd1 vccd1 vccd1 _16855_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout173 _11617_/A2 vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__buf_4
Xfanout184 fanout209/X vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__buf_4
Xfanout195 _12374_/B vssd1 vssd1 vccd1 vccd1 _12377_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ _13873_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _17216_/CLK _15600_/D vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfxtp_1
X_12812_ hold3546/X _12811_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__mux2_1
X_16580_ _18228_/CLK _16580_/D vssd1 vssd1 vccd1 vccd1 _16580_/Q sky130_fd_sc_hd__dfxtp_1
X_13792_ hold4949/X _13880_/B _13791_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ _15531_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__or2_1
X_12743_ hold3035/X _12742_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__mux2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18378_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15462_ _15471_/A _15462_/B _15462_/C _15462_/D vssd1 vssd1 vccd1 vccd1 _15462_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ hold3012/X _12673_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17266_/CLK _17201_/D vssd1 vssd1 vccd1 vccd1 _17201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14413_ _14986_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _14413_/X sky130_fd_sc_hd__or2_1
X_18181_ _18192_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
X_11625_ _12204_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15393_ _15481_/A1 _15385_/X _15392_/X _15481_/B1 _18415_/Q vssd1 vssd1 vccd1 vccd1
+ _15393_/X sky130_fd_sc_hd__a32o_1
X_17132_ _17253_/CLK _17132_/D vssd1 vssd1 vccd1 vccd1 _17132_/Q sky130_fd_sc_hd__dfxtp_1
X_14344_ _14344_/A _14344_/B vssd1 vssd1 vccd1 vccd1 _17971_/D sky130_fd_sc_hd__and2_1
X_11556_ _11652_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ hold4714/X _10073_/B _10506_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10507_/X
+ sky130_fd_sc_hd__o211a_1
X_17063_ _17879_/CLK _17063_/D vssd1 vssd1 vccd1 vccd1 _17063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ hold2080/X _14272_/B _14274_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14275_/X
+ sky130_fd_sc_hd__o211a_1
X_11487_ _12051_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ _18421_/CLK _16014_/D vssd1 vssd1 vccd1 vccd1 _16014_/Q sky130_fd_sc_hd__dfxtp_1
X_13226_ _17579_/Q _17113_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
X_10438_ hold4449/X _10589_/B _10437_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13156_/X hold5900/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
X_10369_ hold5197/X _10628_/B _10368_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _10369_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12204_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__or2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13081_/X _13087_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17529_/D sky130_fd_sc_hd__o21a_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _18025_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
X_12039_ _13392_/A _12039_/B vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__or2_1
X_16916_ _17862_/CLK _16916_/D vssd1 vssd1 vccd1 vccd1 _16916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ _17896_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _18050_/CLK _16847_/D vssd1 vssd1 vccd1 vccd1 _16847_/Q sky130_fd_sc_hd__dfxtp_1
X_16778_ _17981_/CLK _16778_/D vssd1 vssd1 vccd1 vccd1 _16778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15729_ _17669_/CLK _15729_/D vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _12777_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _16236_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _18448_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08201_ _14529_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__or2_1
X_09181_ hold2536/X _09218_/B _09180_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18379_ _18399_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08132_ _15537_/A hold2084/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08063_ hold2805/X _08082_/B _08062_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _08063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3202 _16740_/Q vssd1 vssd1 vccd1 vccd1 hold3202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3213 _13513_/X vssd1 vssd1 vccd1 vccd1 _17624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3224 _11074_/X vssd1 vssd1 vccd1 vccd1 _16848_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3235 _10423_/X vssd1 vssd1 vccd1 vccd1 _16631_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3246 _17470_/Q vssd1 vssd1 vccd1 vccd1 hold3246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2501 _17953_/Q vssd1 vssd1 vccd1 vccd1 hold2501/X sky130_fd_sc_hd__dlygate4sd3_1
X_08965_ hold179/X hold257/X _08965_/S vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__mux2_1
Xhold3257 _17378_/Q vssd1 vssd1 vccd1 vccd1 hold3257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 _09113_/X vssd1 vssd1 vccd1 vccd1 _16171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3268 _11830_/X vssd1 vssd1 vccd1 vccd1 _17100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _08006_/X vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 _15758_/Q vssd1 vssd1 vccd1 vccd1 hold2534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3279 _16745_/Q vssd1 vssd1 vccd1 vccd1 hold3279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 _14037_/X vssd1 vssd1 vccd1 vccd1 _17824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 _09109_/X vssd1 vssd1 vccd1 vccd1 _16169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 _18105_/Q vssd1 vssd1 vccd1 vccd1 hold1811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2556 _08497_/X vssd1 vssd1 vccd1 vccd1 _15877_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07916_ _15539_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07916_/X sky130_fd_sc_hd__or2_1
Xhold1822 _15794_/Q vssd1 vssd1 vccd1 vccd1 hold1822/X sky130_fd_sc_hd__dlygate4sd3_1
X_08896_ hold59/X hold563/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2567 _09300_/X vssd1 vssd1 vccd1 vccd1 _16260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 _07923_/X vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 _17954_/Q vssd1 vssd1 vccd1 vccd1 hold2578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _18095_/Q vssd1 vssd1 vccd1 vccd1 hold1844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 _08255_/X vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1855 _15550_/X vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 _15876_/Q vssd1 vssd1 vccd1 vccd1 hold1866/X sky130_fd_sc_hd__dlygate4sd3_1
X_07847_ _15525_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07847_/X sky130_fd_sc_hd__or2_1
Xhold1877 _15793_/Q vssd1 vssd1 vccd1 vccd1 hold1877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1888 _14591_/X vssd1 vssd1 vccd1 vccd1 _18089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 _18243_/Q vssd1 vssd1 vccd1 vccd1 hold1899/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09517_ hold3177/X _09517_/A2 _09516_/X _15354_/A vssd1 vssd1 vccd1 vccd1 _09517_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09447_/A _09444_/X _09481_/B vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_192_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09379_ _17326_/Q _15479_/A2 _15447_/B1 hold692/X _09378_/X vssd1 vssd1 vccd1 vccd1
+ _09383_/B sky130_fd_sc_hd__a221o_1
X_11410_ hold4397/X _11792_/B _11409_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _12438_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _17288_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ hold4992/X _11726_/B _11340_/X _15506_/A vssd1 vssd1 vccd1 vccd1 _16937_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _15513_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14060_/X sky130_fd_sc_hd__or2_1
X_11272_ hold5633/X _11753_/B _11271_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11272_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5160 _16507_/Q vssd1 vssd1 vccd1 vccd1 hold5160/X sky130_fd_sc_hd__dlygate4sd3_1
X_13011_ hold667/X _13017_/B vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__or2_1
X_10223_ hold1973/X _16565_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__mux2_1
Xhold5171 _16384_/Q vssd1 vssd1 vccd1 vccd1 hold5171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5182 _15383_/X vssd1 vssd1 vccd1 vccd1 _15384_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5193 _16616_/Q vssd1 vssd1 vccd1 vccd1 hold5193/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_70_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4470 _11458_/X vssd1 vssd1 vccd1 vccd1 _16976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4481 _13357_/X vssd1 vssd1 vccd1 vccd1 _17572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10154_ hold2403/X hold3630/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__mux2_1
Xhold4492 _17019_/Q vssd1 vssd1 vccd1 vccd1 hold4492/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3780 _11722_/Y vssd1 vssd1 vccd1 vccd1 _17064_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14962_ _15123_/A _14962_/B vssd1 vssd1 vccd1 vccd1 _14962_/X sky130_fd_sc_hd__or2_1
Xhold3791 _11745_/Y vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17750_ _18461_/CLK hold929/X vssd1 vssd1 vccd1 vccd1 _17750_/Q sky130_fd_sc_hd__dfxtp_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ hold1804/X hold3912/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__mux2_1
X_16701_ _18227_/CLK _16701_/D vssd1 vssd1 vccd1 vccd1 _16701_/Q sky130_fd_sc_hd__dfxtp_1
X_13913_ _13913_/A hold884/X vssd1 vssd1 vccd1 vccd1 hold885/A sky130_fd_sc_hd__and2_1
X_14893_ hold1702/X _14882_/B _14892_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14893_/X
+ sky130_fd_sc_hd__o211a_1
X_17681_ _17745_/CLK _17681_/D vssd1 vssd1 vccd1 vccd1 _17681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _17735_/Q _13844_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__and3_1
X_16632_ _18190_/CLK _16632_/D vssd1 vssd1 vccd1 vccd1 _16632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16563_ _18095_/CLK _16563_/D vssd1 vssd1 vccd1 vccd1 _16563_/Q sky130_fd_sc_hd__dfxtp_1
X_13775_ hold2032/X hold4731/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ hold4159/X _11177_/B _10986_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _10987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18302_ _18422_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_12726_ _12813_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _17418_/D sky130_fd_sc_hd__and2_1
X_15514_ hold2934/X _15560_/A2 _15513_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__o211a_1
X_16494_ _18416_/CLK _16494_/D vssd1 vssd1 vccd1 vccd1 _16494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _15445_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__or2_1
X_18233_ _18233_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _15502_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _17395_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ hold4702/X _11798_/B _11607_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11608_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _17341_/Q _09362_/C _09362_/D hold646/X vssd1 vssd1 vccd1 vccd1 _15376_/X
+ sky130_fd_sc_hd__a22o_1
X_18164_ _18190_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _15506_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _17372_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17115_ _17275_/CLK _17115_/D vssd1 vssd1 vccd1 vccd1 _17115_/Q sky130_fd_sc_hd__dfxtp_1
X_14327_ hold2564/X _14326_/B _14326_/Y _14813_/C1 vssd1 vssd1 vccd1 vccd1 _14327_/X
+ sky130_fd_sc_hd__o211a_1
X_18095_ _18095_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ hold4615/X _11732_/B _11538_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _11539_/X
+ sky130_fd_sc_hd__o211a_1
Xhold407 hold78/X vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__buf_4
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17046_ _17798_/CLK _17046_/D vssd1 vssd1 vccd1 vccd1 _17046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold429 hold572/X vssd1 vssd1 vccd1 vccd1 hold573/A sky130_fd_sc_hd__buf_6
X_14258_ _15099_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13209_ _13209_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__and2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ hold1320/X _14202_/B _14188_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _14189_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 hold799/X vssd1 vssd1 vccd1 vccd1 hold800/A sky130_fd_sc_hd__buf_6
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08750_ _15334_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _15995_/D sky130_fd_sc_hd__and2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _16235_/Q vssd1 vssd1 vccd1 vccd1 hold1107/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _17977_/Q vssd1 vssd1 vccd1 vccd1 hold1118/X sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _18047_/CLK hold625/X vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1129 _08465_/X vssd1 vssd1 vccd1 vccd1 _15861_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08681_ hold126/X hold614/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__mux2_1
X_17879_ _17879_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ hold1112/X _09338_/A2 _09301_/X _12918_/A vssd1 vssd1 vccd1 vccd1 _09302_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _14218_/A hold2540/X _09277_/S vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ _15547_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_160_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08115_ _13905_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09095_ hold1752/X _09106_/B _09094_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _09095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08046_ hold2145/X _08033_/B _08045_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _08046_/X
+ sky130_fd_sc_hd__o211a_1
Xhold930 hold930/A vssd1 vssd1 vccd1 vccd1 hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 hold941/A vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 hold952/A vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3010 _18379_/Q vssd1 vssd1 vccd1 vccd1 hold3010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 hold974/A vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 _12620_/X vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 _12638_/X vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3043 _12935_/X vssd1 vssd1 vccd1 vccd1 _12936_/B sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _11155_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _09997_/Y sky130_fd_sc_hd__nor2_1
Xhold3054 _17452_/Q vssd1 vssd1 vccd1 vccd1 hold3054/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3065 _17456_/Q vssd1 vssd1 vccd1 vccd1 hold3065/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2320 _17830_/Q vssd1 vssd1 vccd1 vccd1 hold2320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2331 _14085_/X vssd1 vssd1 vccd1 vccd1 _17847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3076 _17369_/Q vssd1 vssd1 vccd1 vccd1 hold3076/X sky130_fd_sc_hd__dlygate4sd3_1
X_08948_ _15314_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _16091_/D sky130_fd_sc_hd__and2_1
Xhold3087 _17443_/Q vssd1 vssd1 vccd1 vccd1 hold3087/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2342 _18124_/Q vssd1 vssd1 vccd1 vccd1 hold2342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2353 _08275_/X vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3098 _12977_/X vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2364 _14711_/X vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 _14817_/X vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 _09105_/X vssd1 vssd1 vccd1 vccd1 _16167_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _08402_/X vssd1 vssd1 vccd1 vccd1 _15831_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _18064_/Q vssd1 vssd1 vccd1 vccd1 hold2386/X sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ _12438_/A hold231/X vssd1 vssd1 vccd1 vccd1 _16057_/D sky130_fd_sc_hd__and2_1
Xhold2397 _15665_/Q vssd1 vssd1 vccd1 vccd1 hold2397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 _17912_/Q vssd1 vssd1 vccd1 vccd1 hold1652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1663 _18360_/Q vssd1 vssd1 vccd1 vccd1 hold1663/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _14697_/X vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1685 _15090_/X vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10910_ hold1300/X _16794_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _10911_/B sky130_fd_sc_hd__mux2_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1696 _18094_/Q vssd1 vssd1 vccd1 vccd1 hold1696/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ hold3315/X _12374_/B _11889_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ hold1171/X _16771_/Q _11219_/C vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _13758_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__or2_1
X_10772_ hold1542/X _16748_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_149_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _07809_/X _12510_/Y _13048_/A hold2175/X vssd1 vssd1 vccd1 vccd1 _12511_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ _13779_/A _13491_/B vssd1 vssd1 vccd1 vccd1 _13491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ hold2346/X _15221_/B _15229_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _15230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _12442_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _17314_/D sky130_fd_sc_hd__and2_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15161_ _15215_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _13888_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14112_ hold756/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14112_/X sky130_fd_sc_hd__or2_1
X_11324_ hold1947/X _16932_/Q _11741_/C vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ hold1567/X _15113_/B _15091_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _15092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14043_ hold841/X _14036_/B _14042_/X _13911_/A vssd1 vssd1 vccd1 vccd1 hold842/A
+ sky130_fd_sc_hd__o211a_1
X_11255_ hold2886/X hold3742/X _11735_/C vssd1 vssd1 vccd1 vccd1 _11256_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10206_ _10542_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__or2_1
X_11186_ _16886_/Q _11192_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__and3_1
X_17802_ _17894_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_1
X_10137_ _10548_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__or2_1
X_15994_ _18408_/CLK _15994_/D vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_276_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17887_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17733_ _17739_/CLK _17733_/D vssd1 vssd1 vccd1 vccd1 _17733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _13294_/A _09951_/A _10067_/X vssd1 vssd1 vccd1 vccd1 _10068_/Y sky130_fd_sc_hd__a21oi_1
X_14945_ hold1527/X _14952_/B _14944_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_205_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _17731_/CLK _17664_/D vssd1 vssd1 vccd1 vccd1 _17664_/Q sky130_fd_sc_hd__dfxtp_1
X_14876_ _15215_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14876_/Y sky130_fd_sc_hd__nand2_1
X_16615_ _18214_/CLK _16615_/D vssd1 vssd1 vccd1 vccd1 _16615_/Q sky130_fd_sc_hd__dfxtp_1
X_13827_ hold3651/X _13734_/A _13826_/X vssd1 vssd1 vccd1 vccd1 _13827_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17595_ _17723_/CLK _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16546_ _18220_/CLK _16546_/D vssd1 vssd1 vccd1 vccd1 _16546_/Q sky130_fd_sc_hd__dfxtp_1
X_13758_ _13758_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ hold2841/X hold3519/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16477_ _18358_/CLK _16477_/D vssd1 vssd1 vccd1 vccd1 _16477_/Q sky130_fd_sc_hd__dfxtp_1
X_13689_ _13788_/A _13689_/B vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18216_ _18216_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
X_15428_ hold368/X _09367_/A _15486_/B1 _17346_/Q vssd1 vssd1 vccd1 vccd1 _15428_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18147_ _18215_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
X_15359_ hold306/X _09365_/B _09392_/C hold83/X _15358_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_124_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5907 _17529_/Q vssd1 vssd1 vccd1 vccd1 hold5907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5918 _17535_/Q vssd1 vssd1 vccd1 vccd1 hold5918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5929 _17537_/Q vssd1 vssd1 vccd1 vccd1 hold5929/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _18080_/CLK hold936/X vssd1 vssd1 vccd1 vccd1 hold934/A sky130_fd_sc_hd__dfxtp_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ hold2943/X _16464_/Q _10022_/C vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__mux2_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _17877_/CLK _17029_/D vssd1 vssd1 vccd1 vccd1 _17029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout706 _08970_/A vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__clkbuf_4
X_09851_ hold1410/X _16441_/Q _10001_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__mux2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout717 _14905_/C1 vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__buf_2
Xfanout728 _09011_/A vssd1 vssd1 vccd1 vccd1 _12422_/A sky130_fd_sc_hd__clkbuf_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__buf_4
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _08970_/A hold693/X vssd1 vssd1 vccd1 vccd1 _16020_/D sky130_fd_sc_hd__and2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ hold1486/X _16418_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__mux2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ hold68/X hold401/X _08793_/S vssd1 vssd1 vccd1 vccd1 _08734_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_147_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08730_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _08669_/S sky130_fd_sc_hd__or2_2
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _09063_/A _08595_/B vssd1 vssd1 vccd1 vccd1 _15921_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _15545_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09216_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09147_ hold1907/X _09164_/B _09146_/X _12885_/A vssd1 vssd1 vccd1 vccd1 _09147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09078_ _15519_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _15217_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nand2_1
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 hold771/A vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 hold849/X vssd1 vssd1 vccd1 vccd1 hold850/A sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _11136_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11040_/X sky130_fd_sc_hd__or2_1
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2150 _14781_/X vssd1 vssd1 vccd1 vccd1 _18181_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 _18012_/Q vssd1 vssd1 vccd1 vccd1 hold2161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 _17875_/Q vssd1 vssd1 vccd1 vccd1 hold2172/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _18197_/Q vssd1 vssd1 vccd1 vccd1 hold2183/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ hold2511/X _17508_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _13993_/X vssd1 vssd1 vccd1 vccd1 _17803_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _09318_/X vssd1 vssd1 vccd1 vccd1 _16269_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _15231_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14730_/X sky130_fd_sc_hd__or2_1
X_11942_ hold1740/X hold3427/X _12332_/C vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__mux2_1
Xhold1471 _16255_/Q vssd1 vssd1 vccd1 vccd1 hold1471/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1482 _16160_/Q vssd1 vssd1 vccd1 vccd1 hold1482/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 hold6017/X vssd1 vssd1 vccd1 vccd1 _09447_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ hold1973/X _14664_/B _14660_/Y _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14661_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ hold355/X hold3191/X _12353_/C vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ hold4775/X _13805_/B _13611_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _13612_/X
+ sky130_fd_sc_hd__o211a_1
X_16400_ _18391_/CLK _16400_/D vssd1 vssd1 vccd1 vccd1 _16400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _11031_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__or2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14986_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__or2_1
X_17380_ _17485_/CLK _17380_/D vssd1 vssd1 vccd1 vccd1 _17380_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16331_ _18380_/CLK _16331_/D vssd1 vssd1 vccd1 vccd1 _16331_/Q sky130_fd_sc_hd__dfxtp_1
X_13543_ hold4463/X _13814_/B _13542_/X _09272_/A vssd1 vssd1 vccd1 vccd1 _13543_/X
+ sky130_fd_sc_hd__o211a_1
X_10755_ _11637_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16262_ _17487_/CLK _16262_/D vssd1 vssd1 vccd1 vccd1 _16262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13474_ hold4595/X _13859_/B _13473_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _13474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ _11106_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15213_ _15213_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__or2_1
X_18001_ _18065_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
X_12425_ hold140/X hold710/X _12425_/S vssd1 vssd1 vccd1 vccd1 hold711/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16193_ _17785_/CLK _16193_/D vssd1 vssd1 vccd1 vccd1 _16193_/Q sky130_fd_sc_hd__dfxtp_1
X_15144_ hold1758/X hold609/X _15143_/X _15144_/C1 vssd1 vssd1 vccd1 vccd1 _15144_/X
+ sky130_fd_sc_hd__o211a_1
X_12356_ _17276_/Q _12356_/B _12356_/C vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11688_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or2_1
X_15075_ _15129_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12287_ hold1981/X hold4217/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14026_ _15533_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__or2_1
X_11238_ _12204_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ hold3696/X _11652_/A _11168_/X vssd1 vssd1 vccd1 vccd1 _11169_/Y sky130_fd_sc_hd__a21oi_1
X_15977_ _18423_/CLK _15977_/D vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _17748_/CLK _17716_/D vssd1 vssd1 vccd1 vccd1 _17716_/Q sky130_fd_sc_hd__dfxtp_1
X_14928_ _15197_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _17647_/CLK _17647_/D vssd1 vssd1 vccd1 vccd1 _17647_/Q sky130_fd_sc_hd__dfxtp_1
X_14859_ hold1531/X _14880_/B _14858_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14859_/X
+ sky130_fd_sc_hd__o211a_1
X_08380_ _15549_/A hold1856/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__mux2_1
X_17578_ _17738_/CLK _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16529_ _18268_/CLK _16529_/D vssd1 vssd1 vccd1 vccd1 _16529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09001_ _15454_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _16117_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5704 _11068_/X vssd1 vssd1 vccd1 vccd1 _16846_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5715 _16983_/Q vssd1 vssd1 vccd1 vccd1 hold5715/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5726 _10744_/X vssd1 vssd1 vccd1 vccd1 _16738_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5737 _16949_/Q vssd1 vssd1 vccd1 vccd1 hold5737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5748 _11284_/X vssd1 vssd1 vccd1 vccd1 _16918_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5759 hold5908/X vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__buf_1
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_198_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17827_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09903_ _09903_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__or2_1
Xfanout503 fanout523/X vssd1 vssd1 vccd1 vccd1 _10568_/C sky130_fd_sc_hd__buf_4
Xfanout514 _10601_/C vssd1 vssd1 vccd1 vccd1 _10055_/C sky130_fd_sc_hd__clkbuf_8
Xfanout525 _09340_/X vssd1 vssd1 vccd1 vccd1 _15481_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout536 _09124_/Y vssd1 vssd1 vccd1 vccd1 _09177_/A2 sky130_fd_sc_hd__buf_4
X_09834_ _09948_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_127_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout547 _08443_/B vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__clkbuf_8
Xfanout558 _08217_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__clkbuf_8
Xfanout569 _07990_/B vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__buf_6
XFILLER_0_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09933_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__or2_1
X_08716_ _15364_/A hold155/X vssd1 vssd1 vccd1 vccd1 _15979_/D sky130_fd_sc_hd__and2_1
X_09696_ _09933_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__or2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ hold251/X hold511/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__mux2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ hold149/X hold216/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ hold3967/X _10897_/A2 _10539_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ hold4979/X _10568_/B _10470_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12210_ _12210_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__or2_1
X_13190_ _13190_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__or2_1
X_12141_ _12255_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _13392_/A _12072_/B vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__or2_1
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
X_15900_ _17318_/CLK _15900_/D vssd1 vssd1 vccd1 vccd1 hold524/A sky130_fd_sc_hd__dfxtp_1
X_11023_ hold5538/X _11213_/B _11022_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _11023_/X
+ sky130_fd_sc_hd__o211a_1
X_16880_ _17923_/CLK _16880_/D vssd1 vssd1 vccd1 vccd1 _16880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _17722_/CLK _15831_/D vssd1 vssd1 vccd1 vccd1 _15831_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _17745_/CLK _15762_/D vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfxtp_1
X_12974_ hold3061/X _12973_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__mux2_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 _18382_/Q vssd1 vssd1 vccd1 vccd1 hold1290/X sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ _18013_/CLK _17501_/D vssd1 vssd1 vccd1 vccd1 _17501_/Q sky130_fd_sc_hd__dfxtp_1
X_14713_ hold1212/X _14718_/B _14712_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14713_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _12210_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__or2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _17211_/CLK _15693_/D vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17432_ _17432_/CLK _17432_/D vssd1 vssd1 vccd1 vccd1 _17432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _14984_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__or2_1
X_11856_ _12153_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ hold3938/X _11216_/B _10806_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__o211a_1
X_14575_ hold2785/X _14610_/B _14574_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14575_/X
+ sky130_fd_sc_hd__o211a_1
X_17363_ _17379_/CLK _17363_/D vssd1 vssd1 vccd1 vccd1 _17363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ hold5272/X _12234_/A _11786_/X vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16314_ _16314_/CLK _16314_/D vssd1 vssd1 vccd1 vccd1 _16314_/Q sky130_fd_sc_hd__dfxtp_1
X_13526_ hold2093/X hold4383/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__mux2_1
X_10738_ hold5510/X _11216_/B _10737_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _10738_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17294_ _17329_/CLK _17294_/D vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13457_ hold1114/X _17606_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13458_/B sky130_fd_sc_hd__mux2_1
X_16245_ _17666_/CLK hold237/X vssd1 vssd1 vccd1 vccd1 _16245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10669_ hold3279/X _11156_/B _10668_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _15454_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _17297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ hold875/X hold3822/X _13388_/S vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__mux2_1
X_16176_ _17482_/CLK _16176_/D vssd1 vssd1 vccd1 vccd1 _16176_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput106 hold5879/X vssd1 vssd1 vccd1 vccd1 ki sky130_fd_sc_hd__buf_12
Xoutput117 hold5860/X vssd1 vssd1 vccd1 vccd1 hold5861/A sky130_fd_sc_hd__buf_6
Xoutput128 hold5853/X vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_12
X_12339_ hold5278/X _12051_/A _12338_/X vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__a21oi_1
X_15127_ hold607/X hold656/A vssd1 vssd1 vccd1 vccd1 hold608/A sky130_fd_sc_hd__nor2_1
Xoutput139 _09339_/A vssd1 vssd1 vccd1 vccd1 load_data sky130_fd_sc_hd__buf_12
Xhold3609 _11149_/Y vssd1 vssd1 vccd1 vccd1 _16873_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15058_ _15058_/A hold486/X vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_291_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17253_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2908 _14701_/X vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14009_ hold1625/X _14036_/B _14008_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _14009_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2919 _17758_/Q vssd1 vssd1 vccd1 vccd1 hold2919/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_220_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17893_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07880_ hold1981/X _07865_/B _07879_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _07880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09550_ hold5566/X _10070_/B _09549_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09550_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08501_ hold2088/X _08488_/B _08500_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _08501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09481_ _09482_/B _09481_/B _09481_/C vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_176_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ hold845/X _08433_/B _08431_/Y _08391_/A vssd1 vssd1 vccd1 vccd1 hold846/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08363_ _12810_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _15813_/D sky130_fd_sc_hd__and2_1
XFILLER_0_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ hold1275/X _08336_/A2 _08293_/X _08383_/A vssd1 vssd1 vccd1 vccd1 _08294_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5501 _11278_/X vssd1 vssd1 vccd1 vccd1 _16916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5512 _16486_/Q vssd1 vssd1 vccd1 vccd1 hold5512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5523 _12235_/X vssd1 vssd1 vccd1 vccd1 _17235_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5534 _16853_/Q vssd1 vssd1 vccd1 vccd1 hold5534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4800 _10306_/X vssd1 vssd1 vccd1 vccd1 _16592_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5545 _09901_/X vssd1 vssd1 vccd1 vccd1 _16457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_308_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4811 _17721_/Q vssd1 vssd1 vccd1 vccd1 hold4811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5556 _17142_/Q vssd1 vssd1 vccd1 vccd1 hold5556/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5567 _09550_/X vssd1 vssd1 vccd1 vccd1 _16340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4822 _16742_/Q vssd1 vssd1 vccd1 vccd1 hold4822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4833 _10474_/X vssd1 vssd1 vccd1 vccd1 _16648_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5578 _16496_/Q vssd1 vssd1 vccd1 vccd1 hold5578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4844 _17702_/Q vssd1 vssd1 vccd1 vccd1 hold4844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5589 _09868_/X vssd1 vssd1 vccd1 vccd1 _16446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4855 _11329_/X vssd1 vssd1 vccd1 vccd1 _16933_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4866 _12040_/X vssd1 vssd1 vccd1 vccd1 _17170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout300 _11061_/A vssd1 vssd1 vccd1 vccd1 _11136_/A sky130_fd_sc_hd__buf_4
Xfanout311 fanout337/X vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__clkbuf_4
Xhold4877 _17177_/Q vssd1 vssd1 vccd1 vccd1 hold4877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4888 _11638_/X vssd1 vssd1 vccd1 vccd1 _17036_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout322 _10515_/A vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__buf_4
Xhold4899 _17199_/Q vssd1 vssd1 vccd1 vccd1 hold4899/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout333 fanout337/X vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__clkbuf_4
Xfanout344 _09368_/Y vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__clkbuf_8
Xfanout355 _08669_/S vssd1 vssd1 vccd1 vccd1 _08721_/S sky130_fd_sc_hd__buf_8
Xfanout366 _15149_/B vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__buf_6
X_09817_ hold5458/X _10025_/B _09816_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _09817_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout377 _14962_/B vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__clkbuf_8
Xfanout388 _14734_/Y vssd1 vssd1 vccd1 vccd1 _14772_/B sky130_fd_sc_hd__clkbuf_8
Xfanout399 _14447_/Y vssd1 vssd1 vccd1 vccd1 _14487_/B sky130_fd_sc_hd__buf_6
XFILLER_0_193_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ hold4323/X _10571_/B _09747_/X _15068_/A vssd1 vssd1 vccd1 vccd1 _09748_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ hold3535/X _10601_/B _09678_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09679_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18420_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11710_ hold4815/X _12320_/B _11709_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _17060_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12789_/A _12690_/B vssd1 vssd1 vccd1 vccd1 _17406_/D sky130_fd_sc_hd__and2_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17882_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11641_ hold4613/X _11735_/B _11640_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11641_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14360_/A _14360_/B vssd1 vssd1 vccd1 vccd1 _17979_/D sky130_fd_sc_hd__and2_1
X_11572_ hold5693/X _11762_/B _11571_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _11572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _13311_/A1 _13309_/X _13310_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13311_/X
+ sky130_fd_sc_hd__o211a_1
Xinput19 input19/A vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_10523_ hold2891/X _16665_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__mux2_1
X_14291_ hold1521/X _14333_/A2 _14290_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14291_/X
+ sky130_fd_sc_hd__o211a_1
X_16030_ _18409_/CLK _16030_/D vssd1 vssd1 vccd1 vccd1 _16030_/Q sky130_fd_sc_hd__dfxtp_1
X_13242_ _17581_/Q _17115_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__mux2_1
X_10454_ hold1110/X _16642_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ _13172_/X hold3625/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__mux2_1
X_10385_ hold2419/X _16619_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ hold4935/X _12314_/B _12123_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12124_/X
+ sky130_fd_sc_hd__o211a_1
X_17981_ _17981_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
X_12055_ hold4593/X _12377_/B _12054_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12055_/X
+ sky130_fd_sc_hd__o211a_1
X_16932_ _18427_/CLK _16932_/D vssd1 vssd1 vccd1 vccd1 _16932_/Q sky130_fd_sc_hd__dfxtp_1
X_11006_ hold1195/X _16826_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__mux2_1
X_16863_ _18066_/CLK _16863_/D vssd1 vssd1 vccd1 vccd1 _16863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _17693_/CLK _15814_/D vssd1 vssd1 vccd1 vccd1 _15814_/Q sky130_fd_sc_hd__dfxtp_1
X_16794_ _18061_/CLK _16794_/D vssd1 vssd1 vccd1 vccd1 _16794_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _17708_/CLK _15745_/D vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ _12987_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _17495_/D sky130_fd_sc_hd__and2_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11908_ hold4172/X _13811_/B _11907_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11908_/X
+ sky130_fd_sc_hd__o211a_1
X_15676_ _17908_/CLK _15676_/D vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12918_/A _12888_/B vssd1 vssd1 vccd1 vccd1 _17472_/D sky130_fd_sc_hd__and2_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17419_/CLK _17415_/D vssd1 vssd1 vccd1 vccd1 _17415_/Q sky130_fd_sc_hd__dfxtp_1
X_14627_ _14627_/A hold656/X vssd1 vssd1 vccd1 vccd1 _14668_/B sky130_fd_sc_hd__or2_4
X_18395_ _18395_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ hold5128/X _12356_/B _11838_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _17531_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _17346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _15492_/A _14573_/B hold1801/X vssd1 vssd1 vccd1 vccd1 _14558_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_172_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ _13800_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _17743_/CLK _17277_/D vssd1 vssd1 vccd1 vccd1 _17277_/Q sky130_fd_sc_hd__dfxtp_1
X_14489_ _15169_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14489_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16228_ _18458_/CLK _16228_/D vssd1 vssd1 vccd1 vccd1 _16228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4107 _16945_/Q vssd1 vssd1 vccd1 vccd1 hold4107/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4118 _13510_/X vssd1 vssd1 vccd1 vccd1 _17623_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16159_ _17981_/CLK _16159_/D vssd1 vssd1 vccd1 vccd1 _16159_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4129 _16605_/Q vssd1 vssd1 vccd1 vccd1 hold4129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3406 _17433_/Q vssd1 vssd1 vccd1 vccd1 hold3406/X sky130_fd_sc_hd__dlygate4sd3_1
X_08981_ hold149/X hold199/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__mux2_1
Xhold3417 _13675_/X vssd1 vssd1 vccd1 vccd1 _17678_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3428 _11848_/X vssd1 vssd1 vccd1 vccd1 _17106_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3439 _12533_/X vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2705 _18050_/Q vssd1 vssd1 vccd1 vccd1 hold2705/X sky130_fd_sc_hd__dlygate4sd3_1
X_07932_ hold800/X _07936_/B vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__or2_1
Xhold2716 _14305_/X vssd1 vssd1 vccd1 vccd1 _17952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2727 _15673_/Q vssd1 vssd1 vccd1 vccd1 hold2727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 _18030_/Q vssd1 vssd1 vccd1 vccd1 hold2738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 _15206_/X vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07863_ _15000_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ hold1255/X _16358_/Q _11066_/S vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__mux2_1
X_07794_ _11155_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09533_ _18248_/Q _13150_/A _10028_/C vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09464_ _09463_/A _09461_/X _09481_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _15529_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09395_ _15354_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _16284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08346_ _14850_/A hold1669/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ hold2725/X _08268_/B _08276_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _08277_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6010 _16310_/Q vssd1 vssd1 vccd1 vccd1 hold6010/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6021 _16315_/Q vssd1 vssd1 vccd1 vccd1 hold6021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6032 _16308_/Q vssd1 vssd1 vccd1 vccd1 hold6032/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5320 _11224_/Y vssd1 vssd1 vccd1 vccd1 _16898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_142_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold5331 _16919_/Q vssd1 vssd1 vccd1 vccd1 hold5331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5342 _17043_/Q vssd1 vssd1 vccd1 vccd1 hold5342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5353 _09793_/X vssd1 vssd1 vccd1 vccd1 _16421_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5364 _09532_/X vssd1 vssd1 vccd1 vccd1 _16334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5375 _17171_/Q vssd1 vssd1 vccd1 vccd1 hold5375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4630 _11332_/X vssd1 vssd1 vccd1 vccd1 _16934_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10170_ _10527_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__or2_1
Xhold5386 _09838_/X vssd1 vssd1 vccd1 vccd1 _16436_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4641 _17675_/Q vssd1 vssd1 vccd1 vccd1 hold4641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4652 _13453_/X vssd1 vssd1 vccd1 vccd1 _17604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5397 _17174_/Q vssd1 vssd1 vccd1 vccd1 hold5397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4663 _17039_/Q vssd1 vssd1 vccd1 vccd1 hold4663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4674 _13585_/X vssd1 vssd1 vccd1 vccd1 _17648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3940 _16842_/Q vssd1 vssd1 vccd1 vccd1 hold3940/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4685 _12118_/X vssd1 vssd1 vccd1 vccd1 _17196_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4696 _17196_/Q vssd1 vssd1 vccd1 vccd1 hold4696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3951 _12306_/Y vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3962 _11056_/X vssd1 vssd1 vccd1 vccd1 _16842_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3973 _10408_/X vssd1 vssd1 vccd1 vccd1 _16626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout152 _12911_/S vssd1 vssd1 vccd1 vccd1 _12920_/S sky130_fd_sc_hd__clkbuf_8
Xhold3984 _10780_/X vssd1 vssd1 vccd1 vccd1 _16750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout163 _12302_/B vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__buf_4
Xfanout174 _10852_/A2 vssd1 vssd1 vccd1 vccd1 _11617_/A2 sky130_fd_sc_hd__clkbuf_4
Xhold3995 _16860_/Q vssd1 vssd1 vccd1 vccd1 hold3995/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout185 fanout209/X vssd1 vssd1 vccd1 vccd1 _13868_/B sky130_fd_sc_hd__buf_2
Xfanout196 fanout209/X vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__buf_4
X_13860_ hold4200/X _13764_/A _13859_/X vssd1 vssd1 vccd1 vccd1 _13860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ hold2365/X hold3113/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _13791_/A _13791_/B vssd1 vssd1 vccd1 vccd1 _13791_/X sky130_fd_sc_hd__or2_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ hold1846/X _15560_/A2 _15529_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _15530_/X
+ sky130_fd_sc_hd__o211a_1
X_12742_ _16245_/Q hold3033/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12742_/X sky130_fd_sc_hd__mux2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ hold714/X _09362_/D _09392_/D hold710/X _15460_/X vssd1 vssd1 vccd1 vccd1
+ _15462_/D sky130_fd_sc_hd__a221o_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ hold1854/X _17402_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux2_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17232_/CLK _17200_/D vssd1 vssd1 vccd1 vccd1 _17200_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ hold1627/X hold3433/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__mux2_1
X_14412_ hold5984/X hold209/X hold1054/X _14350_/A vssd1 vssd1 vccd1 vccd1 _14412_/X
+ sky130_fd_sc_hd__o211a_1
X_18180_ _18266_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
X_15392_ _15471_/A _15392_/B _15392_/C _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17131_ _18428_/CLK _17131_/D vssd1 vssd1 vccd1 vccd1 _17131_/Q sky130_fd_sc_hd__dfxtp_1
X_11555_ hold1434/X _17009_/Q _11747_/C vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__mux2_1
X_14343_ hold756/X hold1086/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _10506_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or2_1
X_17062_ _18426_/CLK _17062_/D vssd1 vssd1 vccd1 vccd1 _17062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14274_ _15169_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
X_11486_ hold1079/X hold4001/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_111_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13225_ _13225_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__and2_1
X_16013_ _18423_/CLK _16013_/D vssd1 vssd1 vccd1 vccd1 _16013_/Q sky130_fd_sc_hd__dfxtp_1
X_10437_ _10551_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ hold3696/X _13155_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__mux2_1
X_10368_ _10491_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__or2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ hold2044/X hold4623/X _12299_/C vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13183_/A1 _13085_/X _13086_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _18055_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
X_10299_ _10551_/A _10299_/B vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__or2_1
X_12038_ hold2239/X hold3495/X _13871_/C vssd1 vssd1 vccd1 vccd1 _12039_/B sky130_fd_sc_hd__mux2_1
X_16915_ _17827_/CLK _16915_/D vssd1 vssd1 vccd1 vccd1 _16915_/Q sky130_fd_sc_hd__dfxtp_1
X_17895_ _17895_/CLK hold805/X vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16846_ _18062_/CLK _16846_/D vssd1 vssd1 vccd1 vccd1 _16846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ _18047_/CLK _16777_/D vssd1 vssd1 vccd1 vccd1 _16777_/Q sky130_fd_sc_hd__dfxtp_1
X_13989_ hold760/X _13986_/B _13988_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 hold761/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15728_ _17731_/CLK hold986/X vssd1 vssd1 vccd1 vccd1 hold985/A sky130_fd_sc_hd__dfxtp_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18447_ _18448_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15659_ _17870_/CLK _15659_/D vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfxtp_1
X_08200_ hold2648/X _08213_/B _08199_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08200_/X
+ sky130_fd_sc_hd__o211a_1
X_09180_ _14218_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ _18378_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _08151_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__and2_1
X_17329_ _17329_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 _17329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08062_ _15521_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3203 _10654_/X vssd1 vssd1 vccd1 vccd1 _16708_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3214 _16567_/Q vssd1 vssd1 vccd1 vccd1 hold3214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3225 _17460_/Q vssd1 vssd1 vccd1 vccd1 hold3225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3236 _17359_/Q vssd1 vssd1 vccd1 vccd1 hold3236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3247 _16611_/Q vssd1 vssd1 vccd1 vccd1 hold3247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2502 _14307_/X vssd1 vssd1 vccd1 vccd1 _17953_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08964_ _12420_/A hold344/X vssd1 vssd1 vccd1 vccd1 _16099_/D sky130_fd_sc_hd__and2_1
Xhold2513 _15833_/Q vssd1 vssd1 vccd1 vccd1 hold2513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3258 _17469_/Q vssd1 vssd1 vccd1 vccd1 hold3258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 _18288_/Q vssd1 vssd1 vccd1 vccd1 hold2524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 _17483_/Q vssd1 vssd1 vccd1 vccd1 hold3269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2535 _08247_/X vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07915_ hold2168/X _07918_/B _07914_/X _08149_/A vssd1 vssd1 vccd1 vccd1 _07915_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2546 _15834_/Q vssd1 vssd1 vccd1 vccd1 hold2546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1801 _18074_/Q vssd1 vssd1 vccd1 vccd1 hold1801/X sky130_fd_sc_hd__dlygate4sd3_1
X_08895_ _15374_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _16065_/D sky130_fd_sc_hd__and2_1
Xhold1812 _14623_/X vssd1 vssd1 vccd1 vccd1 _18105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2557 _18438_/Q vssd1 vssd1 vccd1 vccd1 hold2557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _08322_/X vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 _15774_/Q vssd1 vssd1 vccd1 vccd1 hold2568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _15604_/Q vssd1 vssd1 vccd1 vccd1 hold1834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 _14309_/X vssd1 vssd1 vccd1 vccd1 _17954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 _14603_/X vssd1 vssd1 vccd1 vccd1 _18095_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07846_ hold1216/X _07869_/B _07845_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _07846_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1856 _15822_/Q vssd1 vssd1 vccd1 vccd1 hold1856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _08495_/X vssd1 vssd1 vccd1 vccd1 _15876_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1878 _08320_/X vssd1 vssd1 vccd1 vccd1 _15793_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 _17791_/Q vssd1 vssd1 vccd1 vccd1 hold1889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09981_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09447_/A _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09456_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ hold543/X _09367_/A _09386_/D hold715/X vssd1 vssd1 vccd1 vccd1 _09378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_323_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08329_ _15553_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__or2_1
XFILLER_0_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ _11631_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11271_ _12234_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11271_/X sky130_fd_sc_hd__or2_1
Xhold5150 _16419_/Q vssd1 vssd1 vccd1 vccd1 hold5150/X sky130_fd_sc_hd__dlygate4sd3_1
X_13010_ hold1874/X _13003_/Y _13009_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13010_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5161 _09955_/X vssd1 vssd1 vccd1 vccd1 _16475_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10222_ hold4321/X _10589_/B _10221_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10222_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5172 _09586_/X vssd1 vssd1 vccd1 vccd1 _16352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5183 _16512_/Q vssd1 vssd1 vccd1 vccd1 hold5183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5194 _10282_/X vssd1 vssd1 vccd1 vccd1 _16584_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4460 _10228_/X vssd1 vssd1 vccd1 vccd1 _16566_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10153_ hold4240/X _10631_/B _10152_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _10153_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4471 _17742_/Q vssd1 vssd1 vccd1 vccd1 hold4471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4482 _17215_/Q vssd1 vssd1 vccd1 vccd1 hold4482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4493 _11491_/X vssd1 vssd1 vccd1 vccd1 _16987_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3770 _17579_/Q vssd1 vssd1 vccd1 vccd1 hold3770/X sky130_fd_sc_hd__dlygate4sd3_1
X_14961_ hold2473/X _14952_/B _14960_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14961_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3781 _16923_/Q vssd1 vssd1 vccd1 vccd1 hold3781/X sky130_fd_sc_hd__dlygate4sd3_1
X_10084_ hold5148/X _10568_/B _10083_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10084_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3792 _11746_/Y vssd1 vssd1 vccd1 vccd1 _17072_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_4
X_16700_ _18206_/CLK _16700_/D vssd1 vssd1 vccd1 vccd1 _16700_/Q sky130_fd_sc_hd__dfxtp_1
X_13912_ hold883/X _17764_/Q hold244/X vssd1 vssd1 vccd1 vccd1 hold884/A sky130_fd_sc_hd__mux2_1
X_17680_ _17739_/CLK _17680_/D vssd1 vssd1 vccd1 vccd1 _17680_/Q sky130_fd_sc_hd__dfxtp_1
X_14892_ _15123_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14892_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ _18221_/CLK _16631_/D vssd1 vssd1 vccd1 vccd1 _16631_/Q sky130_fd_sc_hd__dfxtp_1
X_13843_ _13873_/A _13843_/B vssd1 vssd1 vccd1 vccd1 _13843_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_187_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16562_ _18210_/CLK _16562_/D vssd1 vssd1 vccd1 vccd1 _16562_/Q sky130_fd_sc_hd__dfxtp_1
X_13774_ hold4993/X _13868_/B _13773_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13774_/X
+ sky130_fd_sc_hd__o211a_1
X_10986_ _11082_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10986_/X sky130_fd_sc_hd__or2_1
X_18301_ _18397_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
X_15513_ _15513_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__or2_1
X_12725_ hold3511/X _12724_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__mux2_1
X_16493_ _18420_/CLK _16493_/D vssd1 vssd1 vccd1 vccd1 _16493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ _18232_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
X_15444_ _15473_/A _15444_/B vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12656_ hold3099/X _12655_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18163_ _18221_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _12153_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__or2_1
X_15375_ hold107/X _15474_/B vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12587_ hold2302/X _12586_/X _12836_/S vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17114_ _17274_/CLK _17114_/D vssd1 vssd1 vccd1 vccd1 _17114_/Q sky130_fd_sc_hd__dfxtp_1
X_14326_ _14774_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _11637_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
X_18094_ _18126_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold408 hold408/A vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold419 hold419/A vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ _17893_/CLK _17045_/D vssd1 vssd1 vccd1 vccd1 _17045_/Q sky130_fd_sc_hd__dfxtp_1
X_11469_ _11667_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__or2_1
X_14257_ hold2844/X _14272_/B _14256_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _14257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _13201_/X _13207_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17544_/D sky130_fd_sc_hd__o21a_1
X_14188_ _15207_/A _14206_/B vssd1 vssd1 vccd1 vccd1 _14188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13138_/X hold3702/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__mux2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _15654_/Q vssd1 vssd1 vccd1 vccd1 hold1108/X sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ _18043_/CLK hold690/X vssd1 vssd1 vccd1 vccd1 hold689/A sky130_fd_sc_hd__dfxtp_1
Xhold1119 _17750_/Q vssd1 vssd1 vccd1 vccd1 hold1119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08680_ _09063_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__and2_1
X_17878_ _17878_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_1
X_16829_ _18032_/CLK _16829_/D vssd1 vssd1 vccd1 vccd1 _16829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09301_ hold949/X _09337_/B vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09232_ hold300/X _15508_/B vssd1 vssd1 vccd1 vccd1 _09232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09163_ hold1923/X _09164_/B _09162_/Y _14360_/A vssd1 vssd1 vccd1 vccd1 _09163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _14854_/A hold2354/X hold196/X vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_160_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09094_ _15535_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08045_ _14786_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__or2_1
Xhold920 hold920/A vssd1 vssd1 vccd1 vccd1 hold920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 hold931/A vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 hold998/X vssd1 vssd1 vccd1 vccd1 hold999/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 la_data_in[7] vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3000 _14585_/X vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3011 _15194_/X vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3022 _17399_/Q vssd1 vssd1 vccd1 vccd1 hold3022/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 _17425_/Q vssd1 vssd1 vccd1 vccd1 hold3033/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3044 _17453_/Q vssd1 vssd1 vccd1 vccd1 hold3044/X sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ _13102_/A _09903_/A _09995_/X vssd1 vssd1 vccd1 vccd1 _09996_/Y sky130_fd_sc_hd__a21oi_1
Xhold2310 _15627_/Q vssd1 vssd1 vccd1 vccd1 hold2310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3055 _17398_/Q vssd1 vssd1 vccd1 vccd1 hold3055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3066 _12839_/X vssd1 vssd1 vccd1 vccd1 _12840_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 _14049_/X vssd1 vssd1 vccd1 vccd1 _17830_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3077 _17422_/Q vssd1 vssd1 vccd1 vccd1 hold3077/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 _16190_/Q vssd1 vssd1 vccd1 vccd1 hold2332/X sky130_fd_sc_hd__dlygate4sd3_1
X_08947_ hold26/X hold598/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__mux2_1
Xhold3088 _12800_/X vssd1 vssd1 vccd1 vccd1 _12801_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2343 _14663_/X vssd1 vssd1 vccd1 vccd1 _18124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3099 _17395_/Q vssd1 vssd1 vccd1 vccd1 hold3099/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2354 _15696_/Q vssd1 vssd1 vccd1 vccd1 hold2354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 _16216_/Q vssd1 vssd1 vccd1 vccd1 hold2365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1620 _09133_/X vssd1 vssd1 vccd1 vccd1 _16179_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2376 _16207_/Q vssd1 vssd1 vccd1 vccd1 hold2376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 hold6021/X vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__buf_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1642 _15883_/Q vssd1 vssd1 vccd1 vccd1 hold1642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 _14536_/X vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ hold32/X _16057_/Q _08932_/S vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__mux2_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 _08051_/X vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1653 _14221_/X vssd1 vssd1 vccd1 vccd1 _17912_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1664 _15154_/X vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1675 _15564_/Q vssd1 vssd1 vccd1 vccd1 hold1675/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _14843_/A hold816/X vssd1 vssd1 vccd1 vccd1 _07829_/Y sky130_fd_sc_hd__nor2_1
Xhold1686 _17846_/Q vssd1 vssd1 vccd1 vccd1 hold1686/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 _14601_/X vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10840_ hold4751/X _11222_/B _10839_/X _14388_/A vssd1 vssd1 vccd1 vccd1 _10840_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ hold5621/X _09992_/B _10770_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _10771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _14556_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12510_/Y sky130_fd_sc_hd__nor2_1
X_13490_ hold1503/X hold4313/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13491_/B sky130_fd_sc_hd__mux2_1
X_12441_ hold14/X hold536/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12442_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15160_ hold1391/X _15161_/B _15159_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15160_/X
+ sky130_fd_sc_hd__o211a_1
X_12372_ hold3828/X _12282_/A _12371_/X vssd1 vssd1 vccd1 vccd1 _12372_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ hold4963/X _12341_/B _11322_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11323_/X
+ sky130_fd_sc_hd__o211a_1
X_14111_ hold1169/X _14148_/B _14110_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _14111_/X
+ sky130_fd_sc_hd__o211a_1
X_15091_ _15199_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15091_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ hold4603/X _11735_/B _11253_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__o211a_1
X_14042_ hold730/X _14050_/B vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__or2_1
X_10205_ hold2187/X _16559_/Q _10637_/C vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ _11218_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__nor2_1
X_17801_ _17892_/CLK hold761/X vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__dfxtp_1
Xhold4290 _11545_/X vssd1 vssd1 vccd1 vccd1 _17005_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10136_ hold1696/X hold3619/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__mux2_1
X_15993_ _18409_/CLK _15993_/D vssd1 vssd1 vccd1 vccd1 _15993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17732_ _17732_/CLK _17732_/D vssd1 vssd1 vccd1 vccd1 _17732_/Q sky130_fd_sc_hd__dfxtp_1
X_10067_ _16513_/Q _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10067_/X sky130_fd_sc_hd__and3_1
X_14944_ _15213_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17663_ _17730_/CLK _17663_/D vssd1 vssd1 vccd1 vccd1 _17663_/Q sky130_fd_sc_hd__dfxtp_1
X_14875_ hold1304/X _14882_/B _14874_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14875_/X
+ sky130_fd_sc_hd__o211a_1
X_16614_ _18204_/CLK _16614_/D vssd1 vssd1 vccd1 vccd1 _16614_/Q sky130_fd_sc_hd__dfxtp_1
X_13826_ _17729_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__and3_1
X_17594_ _17722_/CLK _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_245_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ _18231_/CLK _16545_/D vssd1 vssd1 vccd1 vccd1 _16545_/Q sky130_fd_sc_hd__dfxtp_1
X_13757_ hold1282/X _17706_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__mux2_1
X_10969_ hold5608/X _09992_/B _10968_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _10969_/X
+ sky130_fd_sc_hd__o211a_1
X_12708_ _12777_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _17412_/D sky130_fd_sc_hd__and2_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16476_ _18363_/CLK _16476_/D vssd1 vssd1 vccd1 vccd1 _16476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ hold873/X _17683_/Q _13883_/C vssd1 vssd1 vccd1 vccd1 _13689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ _18215_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15427_ _16095_/Q _09392_/B _09392_/C hold117/X vssd1 vssd1 vccd1 vccd1 _15427_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _12855_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _17389_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _18210_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
X_15358_ hold414/X _09386_/A _15451_/A2 hold698/X vssd1 vssd1 vccd1 vccd1 _15358_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5908 _17545_/Q vssd1 vssd1 vccd1 vccd1 hold5908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5919 _17548_/Q vssd1 vssd1 vccd1 vccd1 hold5919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold205 hold621/X vssd1 vssd1 vccd1 vccd1 hold622/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14309_ hold2578/X _14333_/A2 _14308_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _14309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18077_ _18080_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ hold392/X _15485_/A2 _15447_/B1 _16033_/Q _15288_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 input21/A sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _17844_/CLK _17028_/D vssd1 vssd1 vccd1 vccd1 _17028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout707 _08970_/A vssd1 vssd1 vccd1 vccd1 _12402_/A sky130_fd_sc_hd__clkbuf_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ hold3285/X _11177_/B _09849_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _09850_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 _15172_/C1 vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__buf_4
Xfanout729 _09011_/A vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__clkbuf_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ hold407/X hold692/X _08801_/S vssd1 vssd1 vccd1 vccd1 hold693/A sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ hold5175/X _10067_/B _09780_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09781_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _15454_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _15986_/D sky130_fd_sc_hd__and2_1
X_08663_ _13043_/C _17518_/Q vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_1
XFILLER_0_152_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08594_ hold291/X hold619/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08595_/B sky130_fd_sc_hd__mux2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09215_ hold1830/X _09216_/B _09214_/Y _15534_/C1 vssd1 vssd1 vccd1 vccd1 _09215_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ _15529_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ hold1416/X _09119_/A2 _09076_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _09077_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ hold1901/X _08029_/B _08027_/Y _08139_/A vssd1 vssd1 vccd1 vccd1 _08028_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18460_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold750 la_data_in[10] vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold761 hold761/A vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 hold851/X vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 hold794/A vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ hold5152/X _10073_/B _09978_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09979_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 _14645_/X vssd1 vssd1 vccd1 vccd1 _18115_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2151 _16279_/Q vssd1 vssd1 vccd1 vccd1 hold2151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2162 _14428_/X vssd1 vssd1 vccd1 vccd1 _18012_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2173 _14143_/X vssd1 vssd1 vccd1 vccd1 _17875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12996_/A _12990_/B vssd1 vssd1 vccd1 vccd1 _17506_/D sky130_fd_sc_hd__and2_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2184 _14815_/X vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1450 hold539/X vssd1 vssd1 vccd1 vccd1 input41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2195 _15716_/Q vssd1 vssd1 vccd1 vccd1 hold2195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 _17915_/Q vssd1 vssd1 vccd1 vccd1 hold1461/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ hold4704/X _12323_/B _11940_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11941_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1472 _09290_/X vssd1 vssd1 vccd1 vccd1 _16255_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 _09091_/X vssd1 vssd1 vccd1 vccd1 _16160_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _09407_/X vssd1 vssd1 vccd1 vccd1 _16289_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _15000_/A _14664_/B vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__nand2_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ hold4846/X _12347_/B _11871_/X _12256_/C1 vssd1 vssd1 vccd1 vccd1 _11872_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13611_ _13710_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823_ hold2917/X hold4625/X _11789_/C vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__mux2_1
X_14591_ hold1887/X _14610_/B _14590_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16330_ _18243_/CLK _16330_/D vssd1 vssd1 vccd1 vccd1 _16330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13542_ _13800_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ hold1521/X _16742_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16261_ _17379_/CLK _16261_/D vssd1 vssd1 vccd1 vccd1 _16261_/Q sky130_fd_sc_hd__dfxtp_1
X_13473_ _13764_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__or2_1
X_10685_ hold1144/X hold3604/X _11747_/C vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18000_ _18032_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ hold987/X _15221_/B _15211_/X _15070_/A vssd1 vssd1 vccd1 vccd1 hold988/A
+ sky130_fd_sc_hd__o211a_1
X_12424_ _15284_/A _12424_/B vssd1 vssd1 vccd1 vccd1 _17305_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ _17785_/CLK _16192_/D vssd1 vssd1 vccd1 vccd1 _16192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _15197_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _13822_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__nor2_1
X_11306_ hold351/X hold5272/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__mux2_1
X_12286_ hold4925/X _12314_/B _12285_/X _08137_/A vssd1 vssd1 vccd1 vccd1 _12286_/X
+ sky130_fd_sc_hd__o211a_1
X_15074_ hold207/X hold656/X vssd1 vssd1 vccd1 vccd1 _15123_/B sky130_fd_sc_hd__or2_4
X_11237_ hold1584/X hold3182/X _11717_/C vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__mux2_1
X_14025_ hold1383/X _14040_/B _14024_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14025_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11168_ _11168_/A _11747_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__and3_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ _10548_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__or2_1
X_15976_ _18415_/CLK _15976_/D vssd1 vssd1 vccd1 vccd1 hold530/A sky130_fd_sc_hd__dfxtp_1
X_11099_ hold2754/X hold5050/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17715_ _17715_/CLK _17715_/D vssd1 vssd1 vccd1 vccd1 _17715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14927_ hold1432/X _14946_/B _14926_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _17678_/CLK _17646_/D vssd1 vssd1 vccd1 vccd1 _17646_/Q sky130_fd_sc_hd__dfxtp_1
X_14858_ _15197_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__or2_1
XFILLER_0_187_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13809_ hold3150/X _13713_/A _13808_/X vssd1 vssd1 vccd1 vccd1 _13809_/Y sky130_fd_sc_hd__a21oi_1
X_17577_ _17737_/CLK _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
X_14789_ hold585/X hold655/X vssd1 vssd1 vccd1 vccd1 _14838_/B sky130_fd_sc_hd__or2_4
X_16528_ _18118_/CLK _16528_/D vssd1 vssd1 vccd1 vccd1 _16528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16459_ _18380_/CLK _16459_/D vssd1 vssd1 vccd1 vccd1 _16459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09000_ hold23/X hold676/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18129_ _18225_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5705 _17079_/Q vssd1 vssd1 vccd1 vccd1 hold5705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5716 _11383_/X vssd1 vssd1 vccd1 vccd1 _16951_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5727 _16750_/Q vssd1 vssd1 vccd1 vccd1 hold5727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5738 _11281_/X vssd1 vssd1 vccd1 vccd1 _16917_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5749 _16893_/Q vssd1 vssd1 vccd1 vccd1 hold5749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09902_ hold958/X hold5542/X _09998_/C vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout504 _11093_/S vssd1 vssd1 vccd1 vccd1 _11213_/C sky130_fd_sc_hd__clkbuf_8
Xfanout515 _10601_/C vssd1 vssd1 vccd1 vccd1 _10481_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 _09327_/B vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__clkbuf_4
X_09833_ hold2390/X hold4014/X _10001_/C vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__mux2_1
Xfanout537 _09108_/B vssd1 vssd1 vccd1 vccd1 _09118_/B sky130_fd_sc_hd__clkbuf_4
Xfanout548 _08440_/A2 vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__clkbuf_8
Xfanout559 _08173_/Y vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__buf_6
X_09764_ hold2932/X hold3287/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ hold50/X _15979_/Q _08727_/S vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_167_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18220_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09695_ _18302_/Q hold4293/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__mux2_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _12438_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _15945_/D sky130_fd_sc_hd__and2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _15374_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _15912_/D sky130_fd_sc_hd__and2_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10563_/A _10470_/B vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ hold973/X _09177_/A2 _09128_/X _12855_/A vssd1 vssd1 vccd1 vccd1 hold974/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ hold1126/X _17204_/Q _12332_/C vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ hold1214/X _17181_/Q _13871_/C vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 hold591/A vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _11103_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _17721_/CLK _15830_/D vssd1 vssd1 vccd1 vccd1 _15830_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _17739_/CLK _15761_/D vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfxtp_1
X_12973_ hold2250/X _17502_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux2_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1280 _15863_/Q vssd1 vssd1 vccd1 vccd1 hold1280/X sky130_fd_sc_hd__dlygate4sd3_1
X_17500_ _18013_/CLK _17500_/D vssd1 vssd1 vccd1 vccd1 _17500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 _15200_/X vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ _15213_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14712_/X sky130_fd_sc_hd__or2_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _15672_/Q _17132_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__mux2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _17253_/CLK _15692_/D vssd1 vssd1 vccd1 vccd1 hold919/A sky130_fd_sc_hd__dfxtp_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17432_/CLK _17431_/D vssd1 vssd1 vccd1 vccd1 _17431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ hold1473/X _14664_/B _14642_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14643_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ hold1913/X hold3942/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__mux2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17362_ _17379_/CLK _17362_/D vssd1 vssd1 vccd1 vccd1 _17362_/Q sky130_fd_sc_hd__dfxtp_1
X_10806_ _11121_/A _10806_/B vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__or2_1
X_14574_ _15129_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11786_ _17086_/Q _12329_/B _12329_/C vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16313_ _17503_/CLK _16313_/D vssd1 vssd1 vccd1 vccd1 _16313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ hold4557/X _13805_/B _13524_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _13525_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17293_ _17513_/CLK _17293_/D vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__dfxtp_1
X_10737_ _11121_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__or2_1
X_16244_ _17666_/CLK hold116/X vssd1 vssd1 vccd1 vccd1 _16244_/Q sky130_fd_sc_hd__dfxtp_1
X_13456_ hold5058/X _13856_/B _13455_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13456_/X
+ sky130_fd_sc_hd__o211a_1
X_10668_ _11136_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12407_ hold59/X hold663/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16175_ _18462_/CLK hold803/X vssd1 vssd1 vccd1 vccd1 _16175_/Q sky130_fd_sc_hd__dfxtp_1
X_13387_ hold4498/X _13832_/B _13386_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13387_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10599_ hold3625/X _10548_/A _10598_/X vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__a21oi_1
Xoutput107 hold3989/X vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ hold2381/X _15109_/B _15125_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _15126_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput118 hold3905/X vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_12
Xoutput129 hold3844/X vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_12
X_12338_ _12338_/A _12338_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ hold335/X hold485/X hold302/X vssd1 vssd1 vccd1 vccd1 hold486/A sky130_fd_sc_hd__mux2_1
X_12269_ hold2129/X hold4490/X _13844_/C vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__mux2_1
Xhold2909 _17890_/Q vssd1 vssd1 vccd1 vccd1 hold2909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14008_ _14850_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14008_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_260_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17678_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15959_ _17323_/CLK _15959_/D vssd1 vssd1 vccd1 vccd1 hold451/A sky130_fd_sc_hd__dfxtp_1
X_08500_ _15559_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09480_ hold634/X _09483_/C vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__and2_1
XFILLER_0_187_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ _14950_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17629_ _17629_/CLK _17629_/D vssd1 vssd1 vccd1 vccd1 _17629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ _15531_/A hold1093/X hold122/X vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08293_ _14511_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5502 _16501_/Q vssd1 vssd1 vccd1 vccd1 hold5502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5513 _09892_/X vssd1 vssd1 vccd1 vccd1 _16454_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5524 _16390_/Q vssd1 vssd1 vccd1 vccd1 hold5524/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5535 _10993_/X vssd1 vssd1 vccd1 vccd1 _16821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4801 _17622_/Q vssd1 vssd1 vccd1 vccd1 hold4801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5546 _16764_/Q vssd1 vssd1 vccd1 vccd1 hold5546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4812 _13708_/X vssd1 vssd1 vccd1 vccd1 _17689_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5557 _11860_/X vssd1 vssd1 vccd1 vccd1 _17110_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4823 _10660_/X vssd1 vssd1 vccd1 vccd1 _16710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5568 _16358_/Q vssd1 vssd1 vccd1 vccd1 hold5568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4834 _17000_/Q vssd1 vssd1 vccd1 vccd1 hold4834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5579 _09922_/X vssd1 vssd1 vccd1 vccd1 _16464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4845 _13651_/X vssd1 vssd1 vccd1 vccd1 _17670_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4856 _17160_/Q vssd1 vssd1 vccd1 vccd1 hold4856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4867 hold5814/X vssd1 vssd1 vccd1 vccd1 hold4867/X sky130_fd_sc_hd__clkbuf_4
Xfanout301 _09981_/A vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__buf_4
Xhold4878 _11965_/X vssd1 vssd1 vccd1 vccd1 _17145_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout312 _10557_/A vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__clkbuf_4
Xfanout323 _10515_/A vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__clkbuf_2
Xhold4889 _17657_/Q vssd1 vssd1 vccd1 vccd1 hold4889/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout334 _10422_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__clkbuf_4
Xfanout345 _09368_/Y vssd1 vssd1 vccd1 vccd1 _15471_/A sky130_fd_sc_hd__buf_4
Xfanout356 _08655_/S vssd1 vssd1 vccd1 vccd1 _08661_/S sky130_fd_sc_hd__buf_8
X_09816_ _09924_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__or2_1
Xfanout367 hold608/X vssd1 vssd1 vccd1 vccd1 hold609/A sky130_fd_sc_hd__clkbuf_1
Xfanout378 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__buf_6
Xfanout389 _14724_/B vssd1 vssd1 vccd1 vccd1 _14732_/B sky130_fd_sc_hd__buf_6
X_09747_ _10380_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or2_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _10098_/A _09678_/B vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__or2_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08629_ hold179/X hold418/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__mux2_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11571_ _11667_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11571_/X sky130_fd_sc_hd__or2_1
X_13310_ _13310_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_64_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17313_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ hold4337/X _10646_/B _10521_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14290_ _14970_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13241_ _13241_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10453_ hold4071/X _10643_/B _10452_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13172_ hold5254/X _13171_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
X_10384_ hold4315/X _10558_/A2 _10383_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _10384_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12285_/A _12123_/B vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17980_ _18047_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _12282_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__or2_1
X_16931_ _17907_/CLK _16931_/D vssd1 vssd1 vccd1 vccd1 _16931_/Q sky130_fd_sc_hd__dfxtp_1
X_11005_ hold5050/X _11177_/B _11004_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _11005_/X
+ sky130_fd_sc_hd__o211a_1
X_16862_ _18065_/CLK _16862_/D vssd1 vssd1 vccd1 vccd1 _16862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 hold826/X vssd1 vssd1 vccd1 vccd1 _14854_/A sky130_fd_sc_hd__buf_8
X_15813_ _17723_/CLK _15813_/D vssd1 vssd1 vccd1 vccd1 _15813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16793_ _18208_/CLK _16793_/D vssd1 vssd1 vccd1 vccd1 _16793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _17715_/CLK _15744_/D vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfxtp_1
X_12956_ hold3572/X _12955_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__mux2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18463_ _18463_/A vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _13716_/A _11907_/B vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__or2_1
X_15675_ _17276_/CLK _15675_/D vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ hold3260/X _12886_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12888_/B sky130_fd_sc_hd__mux2_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17414_ _17754_/CLK _17414_/D vssd1 vssd1 vccd1 vccd1 _17414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14627_/A hold655/X vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nor2_1
X_18394_ _18396_/CLK hold979/X vssd1 vssd1 vccd1 vccd1 hold978/A sky130_fd_sc_hd__dfxtp_1
X_11838_ _12267_/A _11838_/B vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 _17345_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14557_ _15492_/A _14573_/B vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11769_ hold5356/X _11694_/A _11768_/X vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ hold2461/X _17623_/Q _13814_/C vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__mux2_1
X_17276_ _17276_/CLK _17276_/D vssd1 vssd1 vccd1 vccd1 _17276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ hold2155/X _14487_/B _14487_/Y _13897_/A vssd1 vssd1 vccd1 vccd1 _14488_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16227_ _18458_/CLK _16227_/D vssd1 vssd1 vccd1 vccd1 _16227_/Q sky130_fd_sc_hd__dfxtp_1
X_13439_ hold2526/X hold3336/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13440_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16158_ _17496_/CLK _16158_/D vssd1 vssd1 vccd1 vccd1 _16158_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4108 _11269_/X vssd1 vssd1 vccd1 vccd1 _16913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4119 _16795_/Q vssd1 vssd1 vccd1 vccd1 hold4119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15109_/A _15109_/B vssd1 vssd1 vccd1 vccd1 _15109_/Y sky130_fd_sc_hd__nand2_1
Xhold3407 _12770_/X vssd1 vssd1 vccd1 vccd1 _12771_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16089_ _17340_/CLK _16089_/D vssd1 vssd1 vccd1 vccd1 hold679/A sky130_fd_sc_hd__dfxtp_1
X_08980_ _15374_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _16107_/D sky130_fd_sc_hd__and2_1
Xhold3418 _17506_/Q vssd1 vssd1 vccd1 vccd1 hold3418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3429 _17489_/Q vssd1 vssd1 vccd1 vccd1 hold3429/X sky130_fd_sc_hd__dlygate4sd3_1
X_07931_ hold2316/X _07924_/B _07930_/X _15502_/A vssd1 vssd1 vccd1 vccd1 _07931_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2706 _14508_/X vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2717 _18033_/Q vssd1 vssd1 vccd1 vccd1 hold2717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 _08067_/X vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2739 _14466_/X vssd1 vssd1 vccd1 vccd1 _18030_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07862_ hold1269/X _07865_/B _07861_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07862_/X
+ sky130_fd_sc_hd__o211a_1
X_09601_ hold4293/X _10022_/B _09600_/X _15038_/A vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ hold5890/X _07788_/A hold1119/X _14556_/A vssd1 vssd1 vccd1 vccd1 _07793_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09532_ hold5363/X _10013_/B _09531_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09463_ _09463_/A _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09472_/D
+ sky130_fd_sc_hd__and4_2
X_08414_ hold2526/X _08440_/A2 _08413_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _08414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ hold5869/A _15481_/B1 _09393_/X _15481_/A1 vssd1 vssd1 vccd1 vccd1 _09394_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _15804_/D sky130_fd_sc_hd__and2_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08276_ hold800/X _08280_/B vssd1 vssd1 vccd1 vccd1 _08276_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6000 _18422_/Q vssd1 vssd1 vccd1 vccd1 hold6000/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6011 _16518_/Q vssd1 vssd1 vccd1 vccd1 hold6011/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6022 _16319_/Q vssd1 vssd1 vccd1 vccd1 hold681/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6033 data_in[4] vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5310 _11202_/Y vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5321 _16927_/Q vssd1 vssd1 vccd1 vccd1 hold5321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5332 _11766_/Y vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5343 _11563_/X vssd1 vssd1 vccd1 vccd1 _17011_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5354 _16429_/Q vssd1 vssd1 vccd1 vccd1 hold5354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4620 _11242_/X vssd1 vssd1 vccd1 vccd1 _16904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5365 _16917_/Q vssd1 vssd1 vccd1 vccd1 hold5365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5376 _11947_/X vssd1 vssd1 vccd1 vccd1 _17139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4631 _17064_/Q vssd1 vssd1 vccd1 vccd1 hold4631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4642 _13570_/X vssd1 vssd1 vccd1 vccd1 _17643_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5387 _16957_/Q vssd1 vssd1 vccd1 vccd1 hold5387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4653 _17205_/Q vssd1 vssd1 vccd1 vccd1 hold4653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5398 _11956_/X vssd1 vssd1 vccd1 vccd1 _17142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4664 _11551_/X vssd1 vssd1 vccd1 vccd1 _17007_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4675 _16593_/Q vssd1 vssd1 vccd1 vccd1 hold4675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3930 _11053_/X vssd1 vssd1 vccd1 vccd1 _16841_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4686 _17029_/Q vssd1 vssd1 vccd1 vccd1 hold4686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3941 _10960_/X vssd1 vssd1 vccd1 vccd1 _16810_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_182_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18228_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4697 _12022_/X vssd1 vssd1 vccd1 vccd1 _17164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3952 _16929_/Q vssd1 vssd1 vccd1 vccd1 hold3952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3963 _17634_/Q vssd1 vssd1 vccd1 vccd1 hold3963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3974 _16752_/Q vssd1 vssd1 vccd1 vccd1 hold3974/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout153 _12911_/S vssd1 vssd1 vccd1 vccd1 _12926_/S sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_111_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18397_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold3985 _16812_/Q vssd1 vssd1 vccd1 vccd1 hold3985/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout164 _09494_/X vssd1 vssd1 vccd1 vccd1 _12302_/B sky130_fd_sc_hd__buf_4
Xhold3996 _11014_/X vssd1 vssd1 vccd1 vccd1 _16828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout175 _10852_/A2 vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__buf_4
Xfanout186 fanout209/X vssd1 vssd1 vccd1 vccd1 _13859_/B sky130_fd_sc_hd__buf_4
Xfanout197 _11783_/B vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__buf_4
X_12810_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _17446_/D sky130_fd_sc_hd__and2_1
X_13790_ hold1859/X hold3539/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13791_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12741_ _12753_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _17423_/D sky130_fd_sc_hd__and2_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15460_ _07805_/A _15477_/A2 _09392_/A hold688/X vssd1 vssd1 vccd1 vccd1 _15460_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12876_/A _12672_/B vssd1 vssd1 vccd1 vccd1 _17400_/D sky130_fd_sc_hd__and2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14411_ _15199_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__or2_1
XFILLER_0_155_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ hold4927/X _12299_/B _11622_/X _08171_/A vssd1 vssd1 vccd1 vccd1 _11623_/X
+ sky130_fd_sc_hd__o211a_1
X_15391_ _16303_/Q _09362_/A _15487_/B1 hold598/X _15390_/X vssd1 vssd1 vccd1 vccd1
+ _15392_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _18445_/CLK _17130_/D vssd1 vssd1 vccd1 vccd1 _17130_/Q sky130_fd_sc_hd__dfxtp_1
X_14342_ _14392_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _17970_/D sky130_fd_sc_hd__and2_1
X_11554_ hold4690/X _11741_/B _11553_/X _14171_/C1 vssd1 vssd1 vccd1 vccd1 _11554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ hold1593/X hold4510/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__mux2_1
X_17061_ _18427_/CLK _17061_/D vssd1 vssd1 vccd1 vccd1 _17061_/Q sky130_fd_sc_hd__dfxtp_1
X_14273_ hold2285/X _14272_/B _14272_/Y _13917_/A vssd1 vssd1 vccd1 vccd1 _14273_/X
+ sky130_fd_sc_hd__o211a_1
X_11485_ hold3890/X _12338_/B _11484_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16012_ _18423_/CLK _16012_/D vssd1 vssd1 vccd1 vccd1 _16012_/Q sky130_fd_sc_hd__dfxtp_1
X_13224_ _13217_/X _13223_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17546_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ hold1292/X _16636_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ _13154_/X _16912_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__mux2_1
X_10367_ hold2901/X hold4779/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ hold4905/X _13811_/B _12105_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _12106_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ hold1212/X _16590_/Q _10589_/C vssd1 vssd1 vccd1 vccd1 _10299_/B sky130_fd_sc_hd__mux2_1
X_13086_ _13086_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__or2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17963_ _18034_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
X_12037_ hold5637/X _12323_/B _12036_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _12037_/X
+ sky130_fd_sc_hd__o211a_1
X_16914_ _17890_/CLK _16914_/D vssd1 vssd1 vccd1 vccd1 _16914_/Q sky130_fd_sc_hd__dfxtp_1
X_17894_ _17894_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_1
X_16845_ _18305_/CLK _16845_/D vssd1 vssd1 vccd1 vccd1 _16845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16776_ _18043_/CLK _16776_/D vssd1 vssd1 vccd1 vccd1 _16776_/Q sky130_fd_sc_hd__dfxtp_1
X_13988_ hold730/X _13992_/B vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _17730_/CLK _15727_/D vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12939_ _12951_/A _12939_/B vssd1 vssd1 vccd1 vccd1 _17489_/D sky130_fd_sc_hd__and2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15658_ _17266_/CLK _15658_/D vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfxtp_1
X_18446_ _18448_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ hold2252/X _14612_/B _14608_/Y _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14609_/X
+ sky130_fd_sc_hd__o211a_1
X_18377_ _18399_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _17205_/CLK _15589_/D vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08130_ _14529_/A hold1603/X _08152_/S vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328_ _18405_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 _17328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08061_ hold2185/X _08082_/B _08060_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _08061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17259_ _18428_/CLK _17259_/D vssd1 vssd1 vccd1 vccd1 _17259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3204 _16654_/Q vssd1 vssd1 vccd1 vccd1 hold3204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3215 _10135_/X vssd1 vssd1 vccd1 vccd1 _16535_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3226 _16343_/Q vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3237 _12548_/X vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08963_ hold71/X _16099_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold344/A sky130_fd_sc_hd__mux2_1
XFILLER_0_110_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3248 _10267_/X vssd1 vssd1 vccd1 vccd1 _16579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2503 _17838_/Q vssd1 vssd1 vccd1 vccd1 hold2503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _08406_/X vssd1 vssd1 vccd1 vccd1 _15833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3259 _17473_/Q vssd1 vssd1 vccd1 vccd1 hold3259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2525 _15005_/X vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2536 _16202_/Q vssd1 vssd1 vccd1 vccd1 hold2536/X sky130_fd_sc_hd__dlygate4sd3_1
X_07914_ _15537_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07914_/X sky130_fd_sc_hd__or2_1
Xhold2547 _08408_/X vssd1 vssd1 vccd1 vccd1 _15834_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1802 _14558_/X vssd1 vssd1 vccd1 vccd1 hold1802/X sky130_fd_sc_hd__dlygate4sd3_1
X_08894_ hold81/X hold716/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__mux2_1
Xhold1813 _18080_/Q vssd1 vssd1 vccd1 vccd1 hold1813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 _15520_/X vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 _15767_/Q vssd1 vssd1 vccd1 vccd1 hold1824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 _08279_/X vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1835 _07921_/X vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07845_ _14517_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07845_/X sky130_fd_sc_hd__or2_1
Xhold1846 _18443_/Q vssd1 vssd1 vccd1 vccd1 hold1846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1857 _18452_/Q vssd1 vssd1 vccd1 vccd1 hold1857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 _17517_/Q vssd1 vssd1 vccd1 vccd1 hold1868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1879 _16221_/Q vssd1 vssd1 vccd1 vccd1 hold1879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09515_ hold956/X _16329_/Q _10763_/S vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ _09444_/X _09446_/B _09481_/B vssd1 vssd1 vccd1 vccd1 _16308_/D sky130_fd_sc_hd__and3b_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ hold5839/A _09342_/B _09342_/Y _09376_/X _12442_/A vssd1 vssd1 vccd1 vccd1
+ _09377_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08328_ hold1271/X _08336_/A2 _08327_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _08328_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ hold873/X _08262_/B _08258_/X _08345_/A vssd1 vssd1 vccd1 vccd1 hold874/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11270_ hold1183/X hold5281/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5140 _16483_/Q vssd1 vssd1 vccd1 vccd1 hold5140/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5151 _09691_/X vssd1 vssd1 vccd1 vccd1 _16387_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10221_ _10551_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5162 _17156_/Q vssd1 vssd1 vccd1 vccd1 hold5162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5173 _17676_/Q vssd1 vssd1 vccd1 vccd1 hold5173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5184 _09970_/X vssd1 vssd1 vccd1 vccd1 _16480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4450 _10438_/X vssd1 vssd1 vccd1 vccd1 _16636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5195 _17644_/Q vssd1 vssd1 vccd1 vccd1 hold5195/X sky130_fd_sc_hd__dlygate4sd3_1
X_10152_ _10542_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or2_1
Xhold4461 hold5816/X vssd1 vssd1 vccd1 vccd1 hold4461/X sky130_fd_sc_hd__clkbuf_4
Xhold4472 _13771_/X vssd1 vssd1 vccd1 vccd1 _17710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4483 _12079_/X vssd1 vssd1 vccd1 vccd1 _17183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4494 _16808_/Q vssd1 vssd1 vccd1 vccd1 hold4494/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3760 _11733_/Y vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__dlygate4sd3_1
X_14960_ _15229_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__or2_1
Xhold3771 _13857_/Y vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__dlygate4sd3_1
X_10083_ _10563_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10083_/X sky130_fd_sc_hd__or2_1
Xhold3782 _11778_/Y vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3793 _17574_/Q vssd1 vssd1 vccd1 vccd1 hold3793/X sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _13911_/A _13911_/B vssd1 vssd1 vccd1 vccd1 _17763_/D sky130_fd_sc_hd__and2_1
X_14891_ hold2570/X _14882_/B _14890_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14891_/X
+ sky130_fd_sc_hd__o211a_1
X_16630_ _18220_/CLK _16630_/D vssd1 vssd1 vccd1 vccd1 _16630_/Q sky130_fd_sc_hd__dfxtp_1
X_13842_ hold3793/X _13764_/A _13841_/X vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16561_ _18215_/CLK _16561_/D vssd1 vssd1 vccd1 vccd1 _16561_/Q sky130_fd_sc_hd__dfxtp_1
X_13773_ _13776_/A _13773_/B vssd1 vssd1 vccd1 vccd1 _13773_/X sky130_fd_sc_hd__or2_1
X_10985_ hold2614/X _16819_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_186_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18300_ _18388_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ hold995/X _15560_/A2 _15511_/X _12885_/A vssd1 vssd1 vccd1 vccd1 hold996/A
+ sky130_fd_sc_hd__o211a_1
X_12724_ hold1081/X hold3486/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16492_ _18334_/CLK _16492_/D vssd1 vssd1 vccd1 vccd1 _16492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18231_ _18231_/CLK hold759/X vssd1 vssd1 vccd1 vccd1 hold758/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15481_/A1 _15435_/X _15442_/X _15490_/B1 _18420_/Q vssd1 vssd1 vccd1 vccd1
+ _15443_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ hold2367/X hold3095/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18162_ _18206_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
X_11606_ _17874_/Q hold4647/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_170_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ hold1894/X _17373_/Q _12679_/S vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17113_ _17583_/CLK _17113_/D vssd1 vssd1 vccd1 vccd1 _17113_/Q sky130_fd_sc_hd__dfxtp_1
X_14325_ hold2423/X _14326_/B _14324_/Y _14344_/A vssd1 vssd1 vccd1 vccd1 _14325_/X
+ sky130_fd_sc_hd__o211a_1
X_18093_ _18229_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ hold2104/X _17003_/Q _11732_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ _17892_/CLK _17044_/D vssd1 vssd1 vccd1 vccd1 _17044_/Q sky130_fd_sc_hd__dfxtp_1
X_14256_ _15205_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__or2_1
X_11468_ hold1132/X _16980_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__mux2_1
X_13207_ _13311_/A1 _13205_/X _13206_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13207_/X
+ sky130_fd_sc_hd__o211a_1
X_10419_ _10515_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__or2_1
X_14187_ hold2824/X _14202_/B _14186_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _14187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11399_ hold1122/X hold5387/X _12338_/C vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__mux2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _17568_/Q _17102_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13138_/X sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13069_ _13068_/X hold3431/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _18043_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1109 _08026_/X vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17877_ _17877_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
X_16828_ _18063_/CLK _16828_/D vssd1 vssd1 vccd1 vccd1 _16828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16759_ _18158_/CLK _16759_/D vssd1 vssd1 vccd1 vccd1 _16759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09300_ hold2566/X _09338_/A2 _09299_/X _12927_/A vssd1 vssd1 vccd1 vccd1 _09300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ hold2205/X _09216_/B _09230_/X _12849_/A vssd1 vssd1 vccd1 vccd1 _09231_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18429_ _18432_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ _15545_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _08139_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__and2_1
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ hold2851/X _09106_/B _09092_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _09093_/X
+ sky130_fd_sc_hd__o211a_1
X_08044_ hold2721/X _08033_/B _08043_/X _12274_/C1 vssd1 vssd1 vccd1 vccd1 _08044_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 hold910/A vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 hold921/A vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold943 hold943/A vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__buf_2
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/A vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3001 _17479_/Q vssd1 vssd1 vccd1 vccd1 hold3001/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold976 hold976/A vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3012 _17401_/Q vssd1 vssd1 vccd1 vccd1 hold3012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 la_data_in[0] vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3023 _17471_/Q vssd1 vssd1 vccd1 vccd1 hold3023/X sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _16489_/Q _09998_/B _09998_/C vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__and3_1
Xhold3034 _12746_/X vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2300 _18169_/Q vssd1 vssd1 vccd1 vccd1 hold2300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3045 _12830_/X vssd1 vssd1 vccd1 vccd1 _12831_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 _07969_/X vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3056 _17406_/Q vssd1 vssd1 vccd1 vccd1 hold3056/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2322 _18182_/Q vssd1 vssd1 vccd1 vccd1 hold2322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08946_ _15374_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _16090_/D sky130_fd_sc_hd__and2_1
Xhold3067 _17459_/Q vssd1 vssd1 vccd1 vccd1 hold3067/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3078 _17385_/Q vssd1 vssd1 vccd1 vccd1 hold3078/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2333 _09155_/X vssd1 vssd1 vccd1 vccd1 _16190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3089 _17404_/Q vssd1 vssd1 vccd1 vccd1 hold3089/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2344 _17910_/Q vssd1 vssd1 vccd1 vccd1 hold2344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 _18328_/Q vssd1 vssd1 vccd1 vccd1 hold1610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2355 _17800_/Q vssd1 vssd1 vccd1 vccd1 hold2355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 _09209_/X vssd1 vssd1 vccd1 vccd1 _16216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 _17836_/Q vssd1 vssd1 vccd1 vccd1 hold1621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 _09423_/X vssd1 vssd1 vccd1 vccd1 _16297_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _15374_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _16056_/D sky130_fd_sc_hd__and2_1
Xhold2377 _09191_/X vssd1 vssd1 vccd1 vccd1 _16207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 _08512_/X vssd1 vssd1 vccd1 vccd1 _15883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 _15612_/Q vssd1 vssd1 vccd1 vccd1 hold2388/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1654 _15642_/Q vssd1 vssd1 vccd1 vccd1 hold1654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2399 _15566_/Q vssd1 vssd1 vccd1 vccd1 hold2399/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1665 _17957_/Q vssd1 vssd1 vccd1 vccd1 hold1665/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1676 _07838_/X vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07828_ _14556_/A hold270/X _14555_/C vssd1 vssd1 vccd1 vccd1 hold815/A sky130_fd_sc_hd__or3_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 _14083_/X vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1698 _18283_/Q vssd1 vssd1 vccd1 vccd1 hold1698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _11067_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _07804_/A _09472_/A _12442_/A _09428_/X vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ _15304_/A _12440_/B vssd1 vssd1 vccd1 vccd1 _17313_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _17281_/Q _12377_/B _12377_/C vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ hold944/X _14160_/B vssd1 vssd1 vccd1 vccd1 _14110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11322_ _12246_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__or2_1
X_15090_ hold1684/X _15113_/B _15089_/X _15026_/A vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14041_ hold2241/X _14040_/B _14040_/Y _14380_/A vssd1 vssd1 vccd1 vccd1 _14041_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _11640_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ hold5032/X _10628_/B _10203_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _10204_/X
+ sky130_fd_sc_hd__o211a_1
X_11184_ hold5251/X _11121_/A _11183_/X vssd1 vssd1 vccd1 vccd1 _11184_/Y sky130_fd_sc_hd__a21oi_1
Xhold4280 _09661_/X vssd1 vssd1 vccd1 vccd1 _16377_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _17903_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_1
X_10135_ hold3214/X _10631_/B _10134_/X _14865_/C1 vssd1 vssd1 vccd1 vccd1 _10135_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4291 _16450_/Q vssd1 vssd1 vccd1 vccd1 hold4291/X sky130_fd_sc_hd__dlygate4sd3_1
X_15992_ _18413_/CLK _15992_/D vssd1 vssd1 vccd1 vccd1 hold597/A sky130_fd_sc_hd__dfxtp_1
Xhold3590 _17365_/Q vssd1 vssd1 vccd1 vccd1 hold3590/X sky130_fd_sc_hd__dlygate4sd3_1
X_14943_ hold831/X _14946_/B _14942_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 hold832/A
+ sky130_fd_sc_hd__o211a_1
X_10066_ _10588_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10066_/Y sky130_fd_sc_hd__nor2_1
X_17731_ _17731_/CLK _17731_/D vssd1 vssd1 vccd1 vccd1 _17731_/Q sky130_fd_sc_hd__dfxtp_1
X_14874_ _15213_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__or2_1
X_17662_ _17694_/CLK _17662_/D vssd1 vssd1 vccd1 vccd1 _17662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16613_ _18235_/CLK _16613_/D vssd1 vssd1 vccd1 vccd1 _16613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13825_ _13864_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nor2_1
X_17593_ _17721_/CLK _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16544_ _18198_/CLK _16544_/D vssd1 vssd1 vccd1 vccd1 _16544_/Q sky130_fd_sc_hd__dfxtp_1
X_13756_ hold5062/X _13880_/B _13755_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _13756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10968_ _11067_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _10968_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ hold3384/X _12706_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__mux2_1
X_16475_ _18396_/CLK _16475_/D vssd1 vssd1 vccd1 vccd1 _16475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13687_ hold5104/X _13880_/B _13686_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13687_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10899_ _11115_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/X sky130_fd_sc_hd__or2_1
X_15426_ _17318_/Q _09357_/A _15446_/B1 hold371/X vssd1 vssd1 vccd1 vccd1 _15426_/X
+ sky130_fd_sc_hd__a22o_1
X_18214_ _18214_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_285_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17844_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12638_ hold3031/X _12637_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18145_ _18388_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
X_15357_ hold462/X _15479_/A2 _09386_/D hold505/X _15356_/X vssd1 vssd1 vccd1 vccd1
+ _15362_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_214_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18032_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12569_ hold3595/X _12568_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5909 _17544_/Q vssd1 vssd1 vccd1 vccd1 hold5909/X sky130_fd_sc_hd__dlygate4sd3_1
X_14308_ _14988_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14308_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18076_ _18080_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
X_15288_ hold217/X _15484_/A2 _15451_/A2 hold309/X vssd1 vssd1 vccd1 vccd1 _15288_/X
+ sky130_fd_sc_hd__a22o_1
Xhold206 hold623/X vssd1 vssd1 vccd1 vccd1 hold624/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17027_ _17904_/CLK _17027_/D vssd1 vssd1 vccd1 vccd1 _17027_/Q sky130_fd_sc_hd__dfxtp_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ hold2699/X _14266_/B _14238_/X _14376_/A vssd1 vssd1 vccd1 vccd1 _14239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 _08970_/A vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout719 _15172_/C1 vssd1 vssd1 vccd1 vccd1 _15036_/A sky130_fd_sc_hd__buf_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _15491_/A hold708/X vssd1 vssd1 vccd1 vccd1 _16019_/D sky130_fd_sc_hd__and2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _10491_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ hold23/X hold631/X _08787_/S vssd1 vssd1 vccd1 vccd1 _08732_/B sky130_fd_sc_hd__mux2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _18059_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
X_08662_ _12426_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _15953_/D sky130_fd_sc_hd__and2_1
XFILLER_0_178_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ _12442_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _15920_/D sky130_fd_sc_hd__and2_1
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _15543_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09145_ hold2542/X _09164_/B _09144_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ _15517_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08027_ _15541_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold740 input49/X vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 hold751/A vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 hold762/A vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold773 hold773/A vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 hold784/A vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__buf_8
Xhold795 hold795/A vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_89_wb_clk_i clkbuf_leaf_90_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17530_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09978_ _10506_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__or2_1
Xhold2130 _07868_/X vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2141 _18131_/Q vssd1 vssd1 vccd1 vccd1 hold2141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08929_ _15304_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _16082_/D sky130_fd_sc_hd__and2_1
Xhold2152 _09338_/X vssd1 vssd1 vccd1 vccd1 _16279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2163 _17832_/Q vssd1 vssd1 vccd1 vccd1 hold2163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2174 hold2209/X vssd1 vssd1 vccd1 vccd1 hold2210/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1440 _18128_/Q vssd1 vssd1 vccd1 vccd1 hold1440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2185 _15670_/Q vssd1 vssd1 vccd1 vccd1 hold2185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 input41/X vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _12036_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__or2_1
Xhold2196 _18321_/Q vssd1 vssd1 vccd1 vccd1 hold2196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1462 _14227_/X vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1473 _18114_/Q vssd1 vssd1 vccd1 vccd1 hold1473/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1484 _15613_/Q vssd1 vssd1 vccd1 vccd1 hold1484/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _18180_/Q vssd1 vssd1 vccd1 vccd1 hold1495/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _12255_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ hold1992/X _17657_/Q _13805_/C vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__mux2_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10822_ hold3922/X _11753_/B _10821_/X _14402_/C1 vssd1 vssd1 vccd1 vccd1 _10822_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14984_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14590_/X sky130_fd_sc_hd__or2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _15819_/Q hold3963/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10753_ hold5480/X _11156_/B _10752_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16260_ _17379_/CLK _16260_/D vssd1 vssd1 vccd1 vccd1 _16260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13472_ _15848_/Q hold3390/X _13859_/C vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__mux2_1
X_10684_ hold5727/X _11201_/B _10683_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ hold735/X _15211_/B vssd1 vssd1 vccd1 vccd1 _15211_/X sky130_fd_sc_hd__or2_1
X_12423_ hold8/X hold151/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12424_/B sky130_fd_sc_hd__mux2_1
X_16191_ _17475_/CLK _16191_/D vssd1 vssd1 vccd1 vccd1 _16191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ hold1410/X _15161_/B _15141_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15142_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12354_ hold3191/X _12285_/A _12353_/X vssd1 vssd1 vccd1 vccd1 _12354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ hold5387/X _12329_/B _11304_/X _14065_/C1 vssd1 vssd1 vccd1 vccd1 _11305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15073_ hold207/X hold656/X vssd1 vssd1 vccd1 vccd1 _15073_/Y sky130_fd_sc_hd__nor2_1
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _15531_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14024_/X sky130_fd_sc_hd__or2_1
X_11236_ hold5036/X _12305_/B _11235_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11236_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _12301_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11167_/Y sky130_fd_sc_hd__nor2_1
X_10118_ hold1597/X hold3625/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__mux2_1
X_15975_ _18413_/CLK _15975_/D vssd1 vssd1 vccd1 vccd1 hold577/A sky130_fd_sc_hd__dfxtp_1
X_11098_ hold4680/X _11192_/B _11097_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _11098_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17714_ _17747_/CLK _17714_/D vssd1 vssd1 vccd1 vccd1 _17714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14926_ _15195_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_1
X_10049_ _16507_/Q _10049_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__and3_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17645_ _17741_/CLK _17645_/D vssd1 vssd1 vccd1 vccd1 _17645_/Q sky130_fd_sc_hd__dfxtp_1
X_14857_ hold1593/X _14880_/B _14856_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14857_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13808_ _17723_/Q _13808_/B _13808_/C vssd1 vssd1 vccd1 vccd1 _13808_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17576_ _17703_/CLK _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
X_14788_ hold585/X hold656/X vssd1 vssd1 vccd1 vccd1 _14788_/Y sky130_fd_sc_hd__nor2_1
X_16527_ _18149_/CLK _16527_/D vssd1 vssd1 vccd1 vccd1 _16527_/Q sky130_fd_sc_hd__dfxtp_1
X_13739_ hold2411/X hold4559/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13740_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16458_ _18371_/CLK _16458_/D vssd1 vssd1 vccd1 vccd1 _16458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15409_ hold450/X _15485_/A2 _15447_/B1 hold328/X _15408_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/C sky130_fd_sc_hd__a221o_1
X_16389_ _18398_/CLK _16389_/D vssd1 vssd1 vccd1 vccd1 _16389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18128_ _18224_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5706 _11671_/X vssd1 vssd1 vccd1 vccd1 _17047_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5717 _16452_/Q vssd1 vssd1 vccd1 vccd1 hold5717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5728 _10684_/X vssd1 vssd1 vccd1 vccd1 _16718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5739 _16952_/Q vssd1 vssd1 vccd1 vccd1 hold5739/X sky130_fd_sc_hd__dlygate4sd3_1
X_18059_ _18059_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09901_ hold5544/X _09998_/B _09900_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout505 _11093_/S vssd1 vssd1 vccd1 vccd1 _11216_/C sky130_fd_sc_hd__clkbuf_8
Xfanout516 fanout523/X vssd1 vssd1 vccd1 vccd1 _10601_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09832_ hold5615/X _10022_/B _09831_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09832_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout527 _09285_/Y vssd1 vssd1 vccd1 vccd1 _09338_/A2 sky130_fd_sc_hd__buf_4
Xfanout538 _09066_/Y vssd1 vssd1 vccd1 vccd1 _09119_/A2 sky130_fd_sc_hd__buf_4
Xfanout549 _08393_/Y vssd1 vssd1 vccd1 vccd1 _08440_/A2 sky130_fd_sc_hd__buf_6
X_09763_ hold5138/X _10049_/B _09762_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09763_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _15491_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _15978_/D sky130_fd_sc_hd__and2_1
X_09694_ hold5681/X _10016_/B _09693_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _09694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ hold149/X hold382/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__mux2_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ hold140/X hold719/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__mux2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_136_wb_clk_i clkbuf_5_26__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18390_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ hold892/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _12426_/A _09059_/B vssd1 vssd1 vccd1 vccd1 _16146_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12070_ hold4439/X _13871_/B _12069_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12070_/X
+ sky130_fd_sc_hd__o211a_1
Xhold570 hold570/A vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 hold581/A vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 hold592/A vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ hold2889/X _16831_/Q _11213_/C vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _17647_/CLK _15760_/D vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _14364_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _17500_/D sky130_fd_sc_hd__and2_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 _07862_/X vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ hold2363/X _14718_/B _14710_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14711_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1281 _08469_/X vssd1 vssd1 vccd1 vccd1 _15863_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ hold5088/X _12305_/B _11922_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11923_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1292 _18194_/Q vssd1 vssd1 vccd1 vccd1 hold1292/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _18426_/CLK _15691_/D vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _15197_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__or2_1
X_17430_ _17432_/CLK _17430_/D vssd1 vssd1 vccd1 vccd1 _17430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ hold3420/X _12362_/B _11853_/X _12142_/C1 vssd1 vssd1 vccd1 vccd1 _11854_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ hold2423/X _16759_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__mux2_1
X_17361_ _17485_/CLK _17361_/D vssd1 vssd1 vccd1 vccd1 _17361_/Q sky130_fd_sc_hd__dfxtp_1
X_14573_ hold281/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14622_/B sky130_fd_sc_hd__nand2_4
X_11785_ _12331_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nor2_1
X_13524_ _13710_/A _13524_/B vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__or2_1
X_16312_ _16314_/CLK _16312_/D vssd1 vssd1 vccd1 vccd1 _16312_/Q sky130_fd_sc_hd__dfxtp_1
X_17292_ _17292_/CLK _17292_/D vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__dfxtp_1
X_10736_ hold1475/X hold5248/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ _17693_/CLK _16243_/D vssd1 vssd1 vccd1 vccd1 hold917/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13455_ _13776_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13455_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ hold1018/X _16713_/Q _10763_/S vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _12420_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _17296_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16174_ _17517_/CLK _16174_/D vssd1 vssd1 vccd1 vccd1 _16174_/Q sky130_fd_sc_hd__dfxtp_1
X_13386_ _13674_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__or2_1
X_10598_ _16690_/Q _10643_/B _10643_/C vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__and3_1
X_15125_ _15233_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__or2_1
Xoutput108 hold5825/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_12
X_12337_ _12343_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12337_/Y sky130_fd_sc_hd__nor2_1
Xoutput119 hold5866/X vssd1 vssd1 vccd1 vccd1 hold5867/A sky130_fd_sc_hd__buf_6
XFILLER_0_142_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15056_ _15056_/A hold303/X vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__and2_1
X_12268_ hold4773/X _12356_/B _12267_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _12268_/X
+ sky130_fd_sc_hd__o211a_1
X_14007_ hold2723/X _14036_/B _14006_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _14007_/X
+ sky130_fd_sc_hd__o211a_1
X_11219_ _16897_/Q _11222_/B _11219_/C vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__and3_1
X_12199_ hold3332/X _12302_/B _12198_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _12199_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput90 _13265_/A vssd1 vssd1 vccd1 vccd1 output90/X sky130_fd_sc_hd__buf_6
XFILLER_0_128_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15958_ _18421_/CLK _15958_/D vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__dfxtp_1
X_14909_ hold956/X hold657/X _14908_/X _15354_/A vssd1 vssd1 vccd1 vccd1 hold957/A
+ sky130_fd_sc_hd__o211a_1
X_15889_ _17345_/CLK _15889_/D vssd1 vssd1 vccd1 vccd1 hold513/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ hold2034/X _08433_/B _08429_/Y _13753_/C1 vssd1 vssd1 vccd1 vccd1 _08430_/X
+ sky130_fd_sc_hd__o211a_1
X_17628_ _17723_/CLK _17628_/D vssd1 vssd1 vccd1 vccd1 _17628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ _12756_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _15812_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17559_ _17719_/CLK _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ hold1638/X _08323_/B _08291_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _08292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5503 _09937_/X vssd1 vssd1 vccd1 vccd1 _16469_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5514 _16499_/Q vssd1 vssd1 vccd1 vccd1 hold5514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5525 _09604_/X vssd1 vssd1 vccd1 vccd1 _16358_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5536 _16858_/Q vssd1 vssd1 vccd1 vccd1 hold5536/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4802 _13411_/X vssd1 vssd1 vccd1 vccd1 _17590_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5547 _10726_/X vssd1 vssd1 vccd1 vccd1 _16732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4813 _17036_/Q vssd1 vssd1 vccd1 vccd1 hold4813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5558 _16868_/Q vssd1 vssd1 vccd1 vccd1 hold5558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4824 _17263_/Q vssd1 vssd1 vccd1 vccd1 hold4824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5569 _09508_/X vssd1 vssd1 vccd1 vccd1 _16326_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4835 _11434_/X vssd1 vssd1 vccd1 vccd1 _16968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4846 _17146_/Q vssd1 vssd1 vccd1 vccd1 hold4846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4857 _11914_/X vssd1 vssd1 vccd1 vccd1 _17128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4868 _15313_/X vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout302 _10779_/A vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4879 _17004_/Q vssd1 vssd1 vccd1 vccd1 hold4879/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout313 _10557_/A vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__clkbuf_4
Xfanout324 fanout337/X vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__buf_2
Xfanout335 _10422_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__buf_4
Xfanout346 _09056_/S vssd1 vssd1 vccd1 vccd1 _09062_/S sky130_fd_sc_hd__buf_8
X_09815_ hold2058/X hold5354/X _10025_/C vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__mux2_1
Xfanout357 _08619_/S vssd1 vssd1 vccd1 vccd1 _08655_/S sky130_fd_sc_hd__buf_8
Xfanout368 hold608/X vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__clkbuf_8
Xfanout379 _14912_/Y vssd1 vssd1 vccd1 vccd1 _14946_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ hold2090/X hold4063/X _10571_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ hold2680/X _16383_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_317_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _15491_/A _08628_/B vssd1 vssd1 vccd1 vccd1 _15936_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _12426_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _15903_/D sky130_fd_sc_hd__and2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ hold1544/X _17014_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13240_ _13233_/X _13239_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_150_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10548_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _13170_/X hold5281/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ _10557_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ hold1548/X hold3400/X _12356_/C vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18072_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12053_ hold2721/X _17175_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__mux2_1
X_16930_ _17905_/CLK _16930_/D vssd1 vssd1 vccd1 vccd1 _16930_/Q sky130_fd_sc_hd__dfxtp_1
X_11004_ _11082_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__or2_1
X_16861_ _18064_/CLK _16861_/D vssd1 vssd1 vccd1 vccd1 _16861_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout880 hold1052/X vssd1 vssd1 vccd1 vccd1 hold1053/A sky130_fd_sc_hd__buf_6
Xfanout891 hold825/X vssd1 vssd1 vccd1 vccd1 hold826/A sky130_fd_sc_hd__clkbuf_2
X_15812_ _17428_/CLK _15812_/D vssd1 vssd1 vccd1 vccd1 _15812_/Q sky130_fd_sc_hd__dfxtp_1
X_16792_ _18061_/CLK _16792_/D vssd1 vssd1 vccd1 vccd1 _16792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _17749_/CLK _15743_/D vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfxtp_1
X_12955_ hold2635/X hold3104/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__mux2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ hold906/X _17126_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__mux2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _18462_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _17262_/CLK _15674_/D vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfxtp_1
X_12886_ hold1742/X hold3259/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__mux2_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17413_ _17754_/CLK _17413_/D vssd1 vssd1 vccd1 vccd1 _17413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11837_ hold941/X hold3825/X _12356_/C vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14625_ hold2218/X _14612_/B _14624_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14625_/X
+ sky130_fd_sc_hd__o211a_1
X_18393_ _18395_/CLK hold931/X vssd1 vssd1 vccd1 vccd1 hold930/A sky130_fd_sc_hd__dfxtp_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17522_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _17344_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14556_/A hold270/X hold241/X vssd1 vssd1 vccd1 vccd1 hold655/A sky130_fd_sc_hd__or3_1
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ _11768_/A _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__and3_1
XFILLER_0_56_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13507_ hold4069/X _13862_/B _13506_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13507_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10719_ _11103_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__or2_1
X_17275_ _17275_/CLK _17275_/D vssd1 vssd1 vccd1 vccd1 _17275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14487_ _15547_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ hold843/X hold4399/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ hold4163/X _13829_/B _13437_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13438_/X
+ sky130_fd_sc_hd__o211a_1
X_16226_ _18458_/CLK _16226_/D vssd1 vssd1 vccd1 vccd1 _16226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16157_ _17506_/CLK _16157_/D vssd1 vssd1 vccd1 vccd1 _16157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ hold4975/X _13847_/B _13368_/X _13753_/C1 vssd1 vssd1 vccd1 vccd1 _13369_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4109 _16626_/Q vssd1 vssd1 vccd1 vccd1 hold4109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ hold2000/X _15109_/B _15107_/Y _15038_/A vssd1 vssd1 vccd1 vccd1 _15108_/X
+ sky130_fd_sc_hd__o211a_1
X_16088_ _17323_/CLK _16088_/D vssd1 vssd1 vccd1 vccd1 hold515/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3408 _16975_/Q vssd1 vssd1 vccd1 vccd1 hold3408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3419 _12989_/X vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07930_ _15553_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__or2_1
X_15039_ _14986_/A hold2263/X hold302/X vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2707 _15637_/Q vssd1 vssd1 vccd1 vccd1 hold2707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 _14472_/X vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2729 _17978_/Q vssd1 vssd1 vccd1 vccd1 hold2729/X sky130_fd_sc_hd__dlygate4sd3_1
X_07861_ _15539_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__or2_1
X_09600_ _09981_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__or2_1
X_07792_ _18460_/Q vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__inv_2
X_09531_ _09933_/A _09531_/B vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _09461_/X _09481_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _16314_/D sky130_fd_sc_hd__and3b_1
X_08413_ _15527_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _07805_/Y _09362_/A _09369_/D _09392_/X vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _14740_/A hold2679/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ hold2352/X _08268_/B _08274_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _08275_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6001 _17524_/Q vssd1 vssd1 vccd1 vccd1 hold6001/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6012 _16316_/Q vssd1 vssd1 vccd1 vccd1 hold6012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6023 data_in[7] vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6034 data_in[8] vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5300 _16739_/Q vssd1 vssd1 vccd1 vccd1 hold5300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5311 _11203_/Y vssd1 vssd1 vccd1 vccd1 _16891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5322 _11790_/Y vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5333 _11767_/Y vssd1 vssd1 vccd1 vccd1 _17079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5344 _17075_/Q vssd1 vssd1 vccd1 vccd1 hold5344/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4610 _10291_/X vssd1 vssd1 vccd1 vccd1 _16587_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5355 _09721_/X vssd1 vssd1 vccd1 vccd1 _16397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4621 _17083_/Q vssd1 vssd1 vccd1 vccd1 hold4621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5366 _11761_/Y vssd1 vssd1 vccd1 vccd1 _17077_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5377 _16500_/Q vssd1 vssd1 vccd1 vccd1 hold5377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4632 _11626_/X vssd1 vssd1 vccd1 vccd1 _17032_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4643 _17260_/Q vssd1 vssd1 vccd1 vccd1 hold4643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5388 _11305_/X vssd1 vssd1 vccd1 vccd1 _16925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5399 _16460_/Q vssd1 vssd1 vccd1 vccd1 hold5399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4654 _12049_/X vssd1 vssd1 vccd1 vccd1 _17173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4665 _16665_/Q vssd1 vssd1 vccd1 vccd1 hold4665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3920 _13851_/Y vssd1 vssd1 vccd1 vccd1 _13852_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4676 _10213_/X vssd1 vssd1 vccd1 vccd1 _16561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3931 _17586_/Q vssd1 vssd1 vccd1 vccd1 hold3931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3942 _17109_/Q vssd1 vssd1 vccd1 vccd1 hold3942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4687 _11521_/X vssd1 vssd1 vccd1 vccd1 _16997_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3953 _11796_/Y vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4698 _16582_/Q vssd1 vssd1 vccd1 vccd1 hold4698/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3964 _13447_/X vssd1 vssd1 vccd1 vccd1 _17602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3975 _10690_/X vssd1 vssd1 vccd1 vccd1 _16720_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout154 _12836_/S vssd1 vssd1 vccd1 vccd1 _12911_/S sky130_fd_sc_hd__buf_4
Xfanout165 _13823_/B vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__buf_4
Xhold3986 _10870_/X vssd1 vssd1 vccd1 vccd1 _16780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3997 _17599_/Q vssd1 vssd1 vccd1 vccd1 hold3997/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout176 _10852_/A2 vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__buf_4
Xfanout187 fanout209/X vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__buf_2
Xfanout198 _11783_/B vssd1 vssd1 vccd1 vccd1 _12338_/B sky130_fd_sc_hd__buf_4
X_09729_ _10779_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_151_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18131_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ hold3038/X _12739_/X _12800_/S vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ hold2864/X _12670_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__mux2_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ hold1294/X hold209/X _14409_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _14410_/X
+ sky130_fd_sc_hd__o211a_1
X_11622_ _12204_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ hold677/X _09367_/A _09392_/A hold568/X vssd1 vssd1 vccd1 vccd1 _15390_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ _15129_/A hold2489/X _14391_/S vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_181_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _12093_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17060_ _17844_/CLK _17060_/D vssd1 vssd1 vccd1 vccd1 _17060_/Q sky130_fd_sc_hd__dfxtp_1
X_10504_ hold4022/X _10646_/B _10503_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o211a_1
X_14272_ _14774_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14272_/Y sky130_fd_sc_hd__nand2_1
X_11484_ _12051_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__or2_1
X_16011_ _16096_/CLK _16011_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13223_ _13311_/A1 _13221_/X _13222_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__o211a_2
X_10435_ hold4236/X _10580_/B _10434_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _10435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13154_ _17570_/Q _17104_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
X_10366_ hold3311/X _11192_/B _10365_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10366_/X
+ sky130_fd_sc_hd__o211a_1
X_12105_ _13716_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__or2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _18158_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
X_13085_ _13084_/X hold3912/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
X_10297_ hold4141/X _10649_/B _10296_/X _14849_/C1 vssd1 vssd1 vccd1 vccd1 _10297_/X
+ sky130_fd_sc_hd__o211a_1
X_12036_ _12036_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__or2_1
X_16913_ _17889_/CLK _16913_/D vssd1 vssd1 vccd1 vccd1 _16913_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_239_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17737_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17893_ _17893_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16844_ _18461_/CLK _16844_/D vssd1 vssd1 vccd1 vccd1 _16844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16775_ _18431_/CLK _16775_/D vssd1 vssd1 vccd1 vccd1 _16775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13987_ hold2355/X _13986_/B _13986_/Y _14191_/C1 vssd1 vssd1 vccd1 vccd1 _13987_/X
+ sky130_fd_sc_hd__o211a_1
X_15726_ _17697_/CLK _15726_/D vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12938_ hold3429/X _12937_/X _13001_/S vssd1 vssd1 vccd1 vccd1 _12938_/X sky130_fd_sc_hd__mux2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18445_ _18445_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15657_ _17902_/CLK _15657_/D vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ hold3330/X _12868_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__mux2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ _15217_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__nand2_1
X_18376_ _18381_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _17268_/CLK _15588_/D vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _18417_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _17327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14539_ _15219_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _15519_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17258_ _18445_/CLK _17258_/D vssd1 vssd1 vccd1 vccd1 _17258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _17448_/CLK _16209_/D vssd1 vssd1 vccd1 vccd1 _16209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17189_ _17221_/CLK _17189_/D vssd1 vssd1 vccd1 vccd1 _17189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3205 _10396_/X vssd1 vssd1 vccd1 vccd1 _16622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3216 _17376_/Q vssd1 vssd1 vccd1 vccd1 hold3216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3227 _10038_/Y vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08962_ _15482_/A hold500/X vssd1 vssd1 vccd1 vccd1 _16098_/D sky130_fd_sc_hd__and2_1
Xhold3238 _16695_/Q vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3249 _17127_/Q vssd1 vssd1 vccd1 vccd1 hold3249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2504 _14067_/X vssd1 vssd1 vccd1 vccd1 _17838_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _17778_/Q vssd1 vssd1 vccd1 vccd1 hold2515/X sky130_fd_sc_hd__dlygate4sd3_1
X_07913_ hold1712/X _07918_/B _07912_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _07913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2526 _15837_/Q vssd1 vssd1 vccd1 vccd1 hold2526/X sky130_fd_sc_hd__dlygate4sd3_1
X_08893_ _12442_/A hold556/X vssd1 vssd1 vccd1 vccd1 _16064_/D sky130_fd_sc_hd__and2_1
Xhold2537 _09181_/X vssd1 vssd1 vccd1 vccd1 _16202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 _18442_/Q vssd1 vssd1 vccd1 vccd1 hold2548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1803 _14559_/X vssd1 vssd1 vccd1 vccd1 _18074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _18244_/Q vssd1 vssd1 vccd1 vccd1 hold2559/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 _14570_/X vssd1 vssd1 vccd1 vccd1 hold1814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1825 _08265_/X vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1836 _18155_/Q vssd1 vssd1 vccd1 vccd1 hold1836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07844_ hold1964/X _07869_/B _07843_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _07844_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1847 _15530_/X vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 _15548_/X vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 _13018_/X vssd1 vssd1 vccd1 vccd1 _17517_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ hold5602/X _09992_/B _09513_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09447_/C _09447_/D _09447_/B vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ hold509/X _15483_/B _09375_/X _18460_/Q vssd1 vssd1 vccd1 vccd1 _09376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ _14330_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ hold735/X _08260_/B vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08189_ _14517_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5130 _17606_/Q vssd1 vssd1 vccd1 vccd1 hold5130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5141 _09883_/X vssd1 vssd1 vccd1 vccd1 _16451_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10220_ hold1191/X hold4165/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__mux2_1
Xhold5152 _16515_/Q vssd1 vssd1 vccd1 vccd1 hold5152/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5163 _11902_/X vssd1 vssd1 vccd1 vccd1 _17124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5174 _13573_/X vssd1 vssd1 vccd1 vccd1 _17644_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5185 hold5815/X vssd1 vssd1 vccd1 vccd1 hold5185/X sky130_fd_sc_hd__clkbuf_4
Xhold4440 _12070_/X vssd1 vssd1 vccd1 vccd1 _17180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10151_ hold2405/X hold3734/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__mux2_1
Xhold5196 _13477_/X vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4451 _16840_/Q vssd1 vssd1 vccd1 vccd1 hold4451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4462 _15303_/X vssd1 vssd1 vccd1 vccd1 _15304_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4473 _16833_/Q vssd1 vssd1 vccd1 vccd1 hold4473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4484 _16484_/Q vssd1 vssd1 vccd1 vccd1 hold4484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3750 _10594_/Y vssd1 vssd1 vccd1 vccd1 _16688_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4495 _10858_/X vssd1 vssd1 vccd1 vccd1 _16776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3761 _11734_/Y vssd1 vssd1 vccd1 vccd1 _17068_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10082_ hold1794/X hold3545/X _10565_/C vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__mux2_1
Xhold3772 _13858_/Y vssd1 vssd1 vccd1 vccd1 _17739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3783 _11779_/Y vssd1 vssd1 vccd1 vccd1 _17083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3794 _13842_/Y vssd1 vssd1 vccd1 vccd1 _13843_/B sky130_fd_sc_hd__dlygate4sd3_1
X_13910_ _15199_/A hold1239/X hold244/X vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__mux2_1
X_14890_ _15229_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14890_/X sky130_fd_sc_hd__or2_1
X_13841_ _17734_/Q _13859_/B _13859_/C vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__and3_1
X_16560_ _18118_/CLK _16560_/D vssd1 vssd1 vccd1 vccd1 _16560_/Q sky130_fd_sc_hd__dfxtp_1
X_13772_ hold2131/X hold4848/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13773_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ hold4228/X _11753_/B _10983_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _10984_/X
+ sky130_fd_sc_hd__o211a_1
X_15511_ hold892/X _15559_/B vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__or2_1
X_12723_ _12813_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _17417_/D sky130_fd_sc_hd__and2_1
X_16491_ _18380_/CLK _16491_/D vssd1 vssd1 vccd1 vccd1 _16491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18230_ _18230_/CLK hold765/X vssd1 vssd1 vccd1 vccd1 hold764/A sky130_fd_sc_hd__dfxtp_1
X_15442_ _15471_/A _15442_/B _15442_/C _15442_/D vssd1 vssd1 vccd1 vccd1 _15442_/X
+ sky130_fd_sc_hd__or4_1
X_12654_ _15502_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _17394_/D sky130_fd_sc_hd__and2_1
XFILLER_0_66_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ hold4399/X _11792_/B _11604_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _11605_/X
+ sky130_fd_sc_hd__o211a_1
X_18161_ _18225_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15373_ _15490_/A1 _15365_/X _15372_/X _15490_/B1 hold5830/A vssd1 vssd1 vccd1 vccd1
+ _15373_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12585_ _12987_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _17371_/D sky130_fd_sc_hd__and2_1
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17112_ _17282_/CLK _17112_/D vssd1 vssd1 vccd1 vccd1 _17112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ hold4339/X _11726_/B _11535_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__o211a_1
X_14324_ _15219_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14324_/Y sky130_fd_sc_hd__nand2_1
X_18092_ _18140_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17043_ _17891_/CLK _17043_/D vssd1 vssd1 vccd1 vccd1 _17043_/Q sky130_fd_sc_hd__dfxtp_1
X_14255_ hold2485/X _14272_/B _14254_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11467_ hold5373/X _11753_/B _11466_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _11467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13206_ _13206_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__or2_1
X_10418_ hold1706/X _16630_/Q _10610_/C vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__mux2_1
X_14186_ _15205_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14186_/X sky130_fd_sc_hd__or2_1
X_11398_ hold4534/X _11741_/B _11397_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _11398_/X
+ sky130_fd_sc_hd__o211a_1
X_13137_ _13137_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__and2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ hold2911/X hold4305/X _10619_/C vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__mux2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _18043_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
X_13068_ hold5590/X _13067_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ hold5015/X _12305_/B _12018_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _12019_/X
+ sky130_fd_sc_hd__o211a_1
X_17876_ _17908_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _18054_/CLK _16827_/D vssd1 vssd1 vccd1 vccd1 _16827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16758_ _18059_/CLK _16758_/D vssd1 vssd1 vccd1 vccd1 _16758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15709_ _17744_/CLK _15709_/D vssd1 vssd1 vccd1 vccd1 hold516/A sky130_fd_sc_hd__dfxtp_1
X_16689_ _18215_/CLK _16689_/D vssd1 vssd1 vccd1 vccd1 _16689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09230_ _15559_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__or2_1
X_18428_ _18428_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09161_ hold1975/X _09164_/B _09160_/Y _14360_/A vssd1 vssd1 vccd1 vccd1 _09161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18359_ _18391_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08112_ _14511_/A hold941/X hold196/X vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _15099_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ _15557_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__or2_1
Xhold900 hold900/A vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 hold911/A vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 hold922/A vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold933 hold933/A vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 hold944/A vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__buf_8
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 input66/X vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 hold977/A vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3002 _12908_/X vssd1 vssd1 vccd1 vccd1 _12909_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3013 _12674_/X vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3024 _12884_/X vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _11155_/A _09994_/B vssd1 vssd1 vccd1 vccd1 _09994_/Y sky130_fd_sc_hd__nor2_1
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3035 _17424_/Q vssd1 vssd1 vccd1 vccd1 hold3035/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2301 _14757_/X vssd1 vssd1 vccd1 vccd1 _18169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3046 _17350_/Q vssd1 vssd1 vccd1 vccd1 hold3046/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2312 _18067_/Q vssd1 vssd1 vccd1 vccd1 hold2312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3057 _17500_/Q vssd1 vssd1 vccd1 vccd1 hold3057/X sky130_fd_sc_hd__dlygate4sd3_1
X_08945_ hold41/X hold535/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__mux2_1
Xhold2323 _14783_/X vssd1 vssd1 vccd1 vccd1 _18182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3068 _12848_/X vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 _15561_/Q vssd1 vssd1 vccd1 vccd1 hold2334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3079 _12626_/X vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1600 _09187_/X vssd1 vssd1 vccd1 vccd1 _16205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2345 _14215_/X vssd1 vssd1 vccd1 vccd1 _17910_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 _15088_/X vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2356 _13987_/X vssd1 vssd1 vccd1 vccd1 _17800_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08876_ hold35/X hold593/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__mux2_1
Xhold2367 _18447_/Q vssd1 vssd1 vccd1 vccd1 hold2367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _14063_/X vssd1 vssd1 vccd1 vccd1 _17836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _15815_/Q vssd1 vssd1 vccd1 vccd1 hold1633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 _16240_/Q vssd1 vssd1 vccd1 vccd1 hold2378/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1644 _15857_/Q vssd1 vssd1 vccd1 vccd1 hold1644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 _07937_/X vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 _08002_/X vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ hold624/A hold279/X hold606/A hold298/X vssd1 vssd1 vccd1 vccd1 _14843_/A
+ sky130_fd_sc_hd__or4b_4
Xhold1666 _14315_/X vssd1 vssd1 vccd1 vccd1 _17957_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1677 _15668_/Q vssd1 vssd1 vccd1 vccd1 hold1677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 _18206_/Q vssd1 vssd1 vccd1 vccd1 hold1688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1699 _14995_/X vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09428_ _09438_/B _16300_/Q vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ hold173/A _15219_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__or3_2
XFILLER_0_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12370_ _13888_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_180_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _17779_/Q hold3871/X _12341_/C vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _14774_/A _14040_/B vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__nand2_1
X_11252_ hold1088/X hold3759/X _11735_/C vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _10491_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _16885_/Q _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__and3_1
Xhold4270 _11548_/X vssd1 vssd1 vccd1 vccd1 _17006_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10134_ _10422_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10134_/X sky130_fd_sc_hd__or2_1
Xhold4281 _17601_/Q vssd1 vssd1 vccd1 vccd1 hold4281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4292 _09784_/X vssd1 vssd1 vccd1 vccd1 _16418_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15991_ _17345_/CLK _15991_/D vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3580 _13558_/X vssd1 vssd1 vccd1 vccd1 _17639_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17730_ _17730_/CLK _17730_/D vssd1 vssd1 vccd1 vccd1 _17730_/Q sky130_fd_sc_hd__dfxtp_1
X_14942_ hold735/X _14962_/B vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or2_1
X_10065_ _13286_/A _10491_/A _10064_/X vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__a21oi_1
Xhold3591 _12566_/X vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__dlygate4sd3_1
X_17661_ _17693_/CLK _17661_/D vssd1 vssd1 vccd1 vccd1 _17661_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2890 _14474_/X vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14873_ hold818/X _14882_/B _14872_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 hold819/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ _18228_/CLK _16612_/D vssd1 vssd1 vccd1 vccd1 _16612_/Q sky130_fd_sc_hd__dfxtp_1
X_13824_ hold3159/X _13737_/A _13823_/X vssd1 vssd1 vccd1 vccd1 _13824_/Y sky130_fd_sc_hd__a21oi_1
X_17592_ _17592_/CLK _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16543_ _18197_/CLK _16543_/D vssd1 vssd1 vccd1 vccd1 _16543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ _13791_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ hold2052/X hold4488/X _11066_/S vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ hold2238/X _17413_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
X_16474_ _18355_/CLK _16474_/D vssd1 vssd1 vccd1 vccd1 _16474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13686_ _13791_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__or2_1
X_10898_ hold2287/X _16790_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _10899_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18213_ _18215_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
X_15425_ _15425_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ hold2443/X _17390_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18144_ _18236_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
X_15356_ _17339_/Q _09362_/C _09362_/D hold534/X vssd1 vssd1 vccd1 vccd1 _15356_/X
+ sky130_fd_sc_hd__a22o_1
X_12568_ hold1648/X hold3107/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11519_ hold2509/X hold4555/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__mux2_1
X_14307_ hold2501/X _14333_/A2 _14306_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _14307_/X
+ sky130_fd_sc_hd__o211a_1
X_18075_ _18080_/CLK hold757/X vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
X_15287_ hold112/X _09357_/A _15484_/B1 hold387/X _15286_/X vssd1 vssd1 vccd1 vccd1
+ _15292_/B sky130_fd_sc_hd__a221o_1
X_12499_ hold65/X _12509_/A2 _12505_/A3 _12498_/X _12426_/A vssd1 vssd1 vccd1 vccd1
+ hold66/A sky130_fd_sc_hd__o311a_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__buf_4
XFILLER_0_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 hold544/X vssd1 vssd1 vccd1 vccd1 hold545/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold31/X vssd1 vssd1 vccd1 vccd1 input31/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17026_ _17905_/CLK _17026_/D vssd1 vssd1 vccd1 vccd1 _17026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14238_ _14972_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_254_wb_clk_i clkbuf_5_17__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17701_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14169_ hold2762/X _14198_/B _14168_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _14169_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 _08970_/A vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__clkbuf_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A _08934_/A vssd1 vssd1 vccd1 vccd1 _08730_/X sky130_fd_sc_hd__or2_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _18190_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08661_ hold291/X hold421/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08662_/B sky130_fd_sc_hd__mux2_1
X_17859_ _17891_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08592_ hold14/X hold523/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ hold1945/X _09216_/B _09212_/Y _15534_/C1 vssd1 vssd1 vccd1 vccd1 _09213_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _15527_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ hold1667/X _09119_/A2 _09074_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08026_ hold1108/X _08029_/B _08025_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _08026_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__buf_4
XFILLER_0_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold730 hold730/A vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold752 input38/X vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 hold763/A vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/A vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 hold796/A vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ hold2756/X hold5140/X _10481_/S vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__mux2_1
Xhold2120 _16253_/Q vssd1 vssd1 vccd1 vccd1 hold2120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2131 _15740_/Q vssd1 vssd1 vccd1 vccd1 hold2131/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2142 _14677_/X vssd1 vssd1 vccd1 vccd1 _18131_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ hold380/X hold633/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__mux2_1
Xhold2153 _15871_/Q vssd1 vssd1 vccd1 vccd1 hold2153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 _14053_/X vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1430 _18260_/Q vssd1 vssd1 vccd1 vccd1 hold1430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2175 hold2211/X vssd1 vssd1 vccd1 vccd1 hold2175/X sky130_fd_sc_hd__clkbuf_2
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1441 _14671_/X vssd1 vssd1 vccd1 vccd1 _18128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2186 _08061_/X vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1452 hold540/X vssd1 vssd1 vccd1 vccd1 hold1452/X sky130_fd_sc_hd__buf_4
Xhold2197 _17825_/Q vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ _15050_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__and2_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1463 _17933_/Q vssd1 vssd1 vccd1 vccd1 hold1463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1474 _14643_/X vssd1 vssd1 vccd1 vccd1 _18114_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _07941_/X vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _14779_/X vssd1 vssd1 vccd1 vccd1 _18180_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ hold1193/X hold3153/X _13388_/S vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_5_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17517_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ _11667_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10821_/X sky130_fd_sc_hd__or2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13540_ hold4385/X _13832_/B _13539_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _13540_/X
+ sky130_fd_sc_hd__o211a_1
X_10752_ _11136_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13471_ hold5179/X _13883_/B _13470_/X _08389_/A vssd1 vssd1 vccd1 vccd1 _13471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _11106_/A _10683_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12422_ _12422_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _17304_/D sky130_fd_sc_hd__and2_1
X_15210_ hold1768/X _15221_/B _15209_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _15210_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16190_ _18432_/CLK _16190_/D vssd1 vssd1 vccd1 vccd1 _16190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15141_ _15195_/A _15149_/B vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__or2_1
X_12353_ _17275_/Q _12356_/B _12353_/C vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11304_ _12234_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11304_/X sky130_fd_sc_hd__or2_1
X_15072_ _15072_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__and2_1
X_12284_ hold2318/X _17252_/Q _13793_/S vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14023_ hold2004/X _14040_/B _14022_/X _14356_/A vssd1 vssd1 vccd1 vccd1 _14023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ _12018_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__or2_1
X_11166_ hold3604/X _11652_/A _11165_/X vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__a21oi_1
X_10117_ hold4407/X _10619_/B _10116_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _10117_/X
+ sky130_fd_sc_hd__o211a_1
X_15974_ _17307_/CLK _15974_/D vssd1 vssd1 vccd1 vccd1 _15974_/Q sky130_fd_sc_hd__dfxtp_1
X_11097_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11097_/X sky130_fd_sc_hd__or2_1
X_17713_ _17745_/CLK _17713_/D vssd1 vssd1 vccd1 vccd1 _17713_/Q sky130_fd_sc_hd__dfxtp_1
X_10048_ _10588_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _16506_/D sky130_fd_sc_hd__nor2_1
X_14925_ hold2983/X _14952_/B _14924_/X _15054_/A vssd1 vssd1 vccd1 vccd1 _14925_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ _17708_/CLK _17644_/D vssd1 vssd1 vccd1 vccd1 _17644_/Q sky130_fd_sc_hd__dfxtp_1
X_14856_ _15195_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13822_/A _13807_/B vssd1 vssd1 vccd1 vccd1 _13807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_188_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _17735_/CLK _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
X_14787_ hold1996/X _14774_/B _14786_/X _14841_/C1 vssd1 vssd1 vccd1 vccd1 _14787_/X
+ sky130_fd_sc_hd__o211a_1
X_11999_ hold2449/X _17157_/Q _13796_/S vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__mux2_1
X_16526_ _18265_/CLK _16526_/D vssd1 vssd1 vccd1 vccd1 _16526_/Q sky130_fd_sc_hd__dfxtp_1
X_13738_ hold4347/X _13832_/B _13737_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13738_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ _18243_/CLK _16457_/D vssd1 vssd1 vccd1 vccd1 _16457_/Q sky130_fd_sc_hd__dfxtp_1
X_13669_ hold5156/X _13859_/B _13668_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ hold325/X _15484_/A2 _15451_/A2 hold474/X vssd1 vssd1 vccd1 vccd1 _15408_/X
+ sky130_fd_sc_hd__a22o_1
X_16388_ _18397_/CLK _16388_/D vssd1 vssd1 vccd1 vccd1 _16388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18127_ _18183_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15339_ hold577/X _15485_/A2 _15447_/B1 hold718/X _15338_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/C sky130_fd_sc_hd__a221o_1
Xhold5707 _17014_/Q vssd1 vssd1 vccd1 vccd1 hold5707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5718 _09790_/X vssd1 vssd1 vccd1 vccd1 _16420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5729 _17015_/Q vssd1 vssd1 vccd1 vccd1 hold5729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058_ _18067_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09900_ _09903_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__or2_1
X_17009_ _17889_/CLK _17009_/D vssd1 vssd1 vccd1 vccd1 _17009_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout506 _10610_/C vssd1 vssd1 vccd1 vccd1 _11093_/S sky130_fd_sc_hd__buf_4
Xfanout517 _10649_/C vssd1 vssd1 vccd1 vccd1 _10589_/C sky130_fd_sc_hd__clkbuf_8
X_09831_ _09987_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__or2_1
Xfanout528 _09285_/Y vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__buf_4
Xfanout539 _09066_/Y vssd1 vssd1 vccd1 vccd1 _09106_/B sky130_fd_sc_hd__buf_4
XFILLER_0_158_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09762_ _09954_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__or2_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ hold251/X hold590/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__mux2_1
X_09693_ _09987_/A _09693_/B vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08644_ _15314_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _15944_/D sky130_fd_sc_hd__and2_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08575_ _15334_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _15911_/D sky130_fd_sc_hd__and2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_176_wb_clk_i clkbuf_5_29__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18003_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ hold2530/X _09177_/A2 _09126_/X _12855_/A vssd1 vssd1 vccd1 vccd1 _09127_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_105_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17314_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09058_ hold380/X hold642/X _09062_/S vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ hold949/X _08045_/B vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__or2_1
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold571 hold571/A vssd1 vssd1 vccd1 vccd1 input50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 hold582/A vssd1 vssd1 vccd1 vccd1 input56/A sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ hold5478/X _11762_/B _11019_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o211a_1
Xhold593 hold593/A vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ hold3057/X _12970_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12971_/X sky130_fd_sc_hd__mux2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 hold1260/A vssd1 vssd1 vccd1 vccd1 input40/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _15103_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14710_/X sky130_fd_sc_hd__or2_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1271 _15797_/Q vssd1 vssd1 vccd1 vccd1 hold1271/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _15735_/Q vssd1 vssd1 vccd1 vccd1 hold1282/X sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _12018_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__or2_1
Xhold1293 _14809_/X vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _17170_/CLK _15690_/D vssd1 vssd1 vccd1 vccd1 _15690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641_ hold2476/X _14664_/B _14640_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _14641_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _12243_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17360_ _17485_/CLK _17360_/D vssd1 vssd1 vccd1 vccd1 _17360_/Q sky130_fd_sc_hd__dfxtp_1
X_10804_ hold4791/X _11192_/B _10803_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _10804_/X
+ sky130_fd_sc_hd__o211a_1
X_11784_ hold3613/X _12234_/A _11783_/X vssd1 vssd1 vccd1 vccd1 _11784_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ hold281/X _14573_/B vssd1 vssd1 vccd1 vccd1 _14572_/X sky130_fd_sc_hd__and2_1
XFILLER_0_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16311_ _16314_/CLK _16311_/D vssd1 vssd1 vccd1 vccd1 _16311_/Q sky130_fd_sc_hd__dfxtp_1
X_13523_ hold1093/X _17628_/Q _13805_/C vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__mux2_1
X_17291_ _18406_/CLK _17291_/D vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__dfxtp_1
X_10735_ hold5452/X _11213_/B _10734_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _10735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _17428_/CLK _16242_/D vssd1 vssd1 vccd1 vccd1 _16242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ hold833/X hold4783/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__mux2_1
X_10666_ hold4547/X _10852_/A2 _10665_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _10666_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ hold81/X hold698/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__mux2_1
X_13385_ hold2153/X hold3814/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__mux2_1
X_16173_ _17516_/CLK _16173_/D vssd1 vssd1 vccd1 vccd1 _16173_/Q sky130_fd_sc_hd__dfxtp_1
X_10597_ _10651_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10597_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ hold1332/X _15113_/B _15123_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _15124_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput109 hold5185/X vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12336_ hold3942/X _12246_/A _12335_/X vssd1 vssd1 vccd1 vccd1 _12336_/Y sky130_fd_sc_hd__a21oi_1
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12267_/X sky130_fd_sc_hd__or2_1
X_15055_ hold235/X _18313_/Q hold302/A vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__mux2_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14006_ _14740_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__or2_1
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__nor2_1
X_12198_ _12210_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__or2_1
Xoutput80 _13193_/A vssd1 vssd1 vccd1 vccd1 output80/X sky130_fd_sc_hd__buf_6
Xoutput91 _13273_/A vssd1 vssd1 vccd1 vccd1 output91/X sky130_fd_sc_hd__buf_6
X_11149_ _11155_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ _17302_/CLK _15957_/D vssd1 vssd1 vccd1 vccd1 _15957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14908_ hold826/X _14910_/B vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__or2_1
X_15888_ _17345_/CLK _15888_/D vssd1 vssd1 vccd1 vccd1 hold509/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17627_ _17691_/CLK _17627_/D vssd1 vssd1 vccd1 vccd1 _17627_/Q sky130_fd_sc_hd__dfxtp_1
X_14839_ hold1337/X _14822_/B _14838_/X _14857_/C1 vssd1 vssd1 vccd1 vccd1 _14839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08360_ _15529_/A hold1843/X hold122/X vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__mux2_1
X_17558_ _17718_/CLK _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16509_ _18358_/CLK _16509_/D vssd1 vssd1 vccd1 vccd1 _16509_/Q sky130_fd_sc_hd__dfxtp_1
X_08291_ _14850_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17489_ _17517_/CLK _17489_/D vssd1 vssd1 vccd1 vccd1 _17489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5504 _17042_/Q vssd1 vssd1 vccd1 vccd1 hold5504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5515 _09931_/X vssd1 vssd1 vccd1 vccd1 _16467_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5526 _16832_/Q vssd1 vssd1 vccd1 vccd1 hold5526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5537 _11008_/X vssd1 vssd1 vccd1 vccd1 _16826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4803 _17168_/Q vssd1 vssd1 vccd1 vccd1 hold4803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5548 _16811_/Q vssd1 vssd1 vccd1 vccd1 hold5548/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4814 _11542_/X vssd1 vssd1 vccd1 vccd1 _17004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5559 _11038_/X vssd1 vssd1 vccd1 vccd1 _16836_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4825 _12223_/X vssd1 vssd1 vccd1 vccd1 _17231_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4836 _17625_/Q vssd1 vssd1 vccd1 vccd1 hold4836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4847 _11872_/X vssd1 vssd1 vccd1 vccd1 _17114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4858 _16581_/Q vssd1 vssd1 vccd1 vccd1 hold4858/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4869 _17217_/Q vssd1 vssd1 vccd1 vccd1 hold4869/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout303 _10779_/A vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__buf_4
Xfanout314 fanout337/X vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__buf_2
Xfanout325 _09951_/A vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__clkbuf_4
Xfanout336 fanout337/X vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__clkbuf_4
Xfanout347 _09028_/S vssd1 vssd1 vccd1 vccd1 _09056_/S sky130_fd_sc_hd__buf_8
X_09814_ hold5399/X _10013_/B _09813_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09814_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout358 _08590_/S vssd1 vssd1 vccd1 vccd1 _08594_/S sky130_fd_sc_hd__buf_8
Xfanout369 _15123_/B vssd1 vssd1 vccd1 vccd1 _15125_/B sky130_fd_sc_hd__clkbuf_8
X_09745_ hold5350/X _10013_/B _09744_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09745_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ hold3328/X _11177_/B _09675_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08627_ hold71/X hold543/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08628_/B sky130_fd_sc_hd__mux2_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ hold59/X hold709/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ hold2279/X _08488_/B _08488_/Y _08143_/A vssd1 vssd1 vccd1 vccd1 _08489_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ hold1555/X hold3924/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ hold2226/X hold4016/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _17572_/Q _17106_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__mux2_1
X_10382_ hold2668/X hold3558/X _11177_/C vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ hold5034/X _12311_/B _12120_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__o211a_1
X_12052_ hold5564/X _12338_/B _12051_/X _13925_/A vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o211a_1
Xhold390 hold390/A vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ hold2971/X _16825_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _18063_/CLK _16860_/D vssd1 vssd1 vccd1 vccd1 _16860_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout870 _07781_/Y vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__buf_12
X_15811_ _17725_/CLK _15811_/D vssd1 vssd1 vccd1 vccd1 _15811_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout881 hold967/X vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__buf_8
Xfanout892 hold490/X vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__buf_8
X_16791_ _18158_/CLK _16791_/D vssd1 vssd1 vccd1 vccd1 _16791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _17745_/CLK _15742_/D vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12996_/A _12954_/B vssd1 vssd1 vccd1 vccd1 _17494_/D sky130_fd_sc_hd__and2_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1090 _13006_/X vssd1 vssd1 vccd1 vccd1 _17511_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ hold4637/X _12308_/B _11904_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__o211a_1
X_18461_ _18461_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _17232_/CLK _15673_/D vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12885_/A _12885_/B vssd1 vssd1 vccd1 vccd1 _17471_/D sky130_fd_sc_hd__and2_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17412_ _17435_/CLK _17412_/D vssd1 vssd1 vccd1 vccd1 _17412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14786_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__or2_1
X_18392_ _18392_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11836_ hold3404/X _12356_/B _11835_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _11836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17343_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 _17343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _18461_/Q _14555_/B _14555_/C vssd1 vssd1 vccd1 vccd1 _14573_/B sky130_fd_sc_hd__and3_4
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11791_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _13767_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__or2_1
X_17274_ _17274_/CLK _17274_/D vssd1 vssd1 vccd1 vccd1 _17274_/Q sky130_fd_sc_hd__dfxtp_1
X_10718_ hold1463/X hold5297/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__mux2_1
X_14486_ hold2350/X _14487_/B _14485_/Y _14907_/C1 vssd1 vssd1 vccd1 vccd1 _14486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11698_ hold4409/X _12341_/B _11697_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11698_/X
+ sky130_fd_sc_hd__o211a_1
X_16225_ _17456_/CLK _16225_/D vssd1 vssd1 vccd1 vccd1 _16225_/Q sky130_fd_sc_hd__dfxtp_1
X_13437_ _13734_/A _13437_/B vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _16707_/Q _10649_/B _10649_/C vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__and3_1
XFILLER_0_130_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16156_ _17506_/CLK _16156_/D vssd1 vssd1 vccd1 vccd1 _16156_/Q sky130_fd_sc_hd__dfxtp_1
X_13368_ _13758_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__or2_1
X_15107_ _15541_/A _15109_/B vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__nand2_1
X_12319_ _13822_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__nor2_1
X_16087_ _17314_/CLK _16087_/D vssd1 vssd1 vccd1 vccd1 hold612/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13299_ _13298_/X hold5903/X _13307_/S vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__mux2_1
Xhold3409 _11359_/X vssd1 vssd1 vccd1 vccd1 _16943_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15038_ _15038_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2708 _07989_/X vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2719 _18278_/Q vssd1 vssd1 vccd1 vccd1 hold2719/X sky130_fd_sc_hd__dlygate4sd3_1
X_07860_ hold2291/X _07865_/B _07859_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07860_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07791_ hold241/X vssd1 vssd1 vccd1 vccd1 _14555_/C sky130_fd_sc_hd__inv_2
XFILLER_0_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16989_ _17891_/CLK _16989_/D vssd1 vssd1 vccd1 vccd1 _16989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09530_ hold2923/X _13142_/A _10010_/C vssd1 vssd1 vccd1 vccd1 _09531_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_155_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__and3_1
X_08412_ hold2562/X _08440_/A2 _08411_/X _08373_/A vssd1 vssd1 vccd1 vccd1 _08412_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ _09392_/A _09392_/B _09392_/C _09392_/D vssd1 vssd1 vccd1 vccd1 _09392_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_47_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08343_ _08345_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08274_ _15553_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6002 becStatus[0] vssd1 vssd1 vccd1 vccd1 hold6002/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6013 data_in[0] vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6024 data_in[24] vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6035 _16306_/Q vssd1 vssd1 vccd1 vccd1 hold6035/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5301 _11226_/Y vssd1 vssd1 vccd1 vccd1 _11227_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5312 _16718_/Q vssd1 vssd1 vccd1 vccd1 hold5312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5323 _11791_/Y vssd1 vssd1 vccd1 vccd1 _17087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5334 _17021_/Q vssd1 vssd1 vccd1 vccd1 hold5334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4600 _11974_/X vssd1 vssd1 vccd1 vccd1 _17148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5345 _11659_/X vssd1 vssd1 vccd1 vccd1 _17043_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5356 _16920_/Q vssd1 vssd1 vccd1 vccd1 hold5356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4611 _16971_/Q vssd1 vssd1 vccd1 vccd1 hold4611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4622 _11683_/X vssd1 vssd1 vccd1 vccd1 _17051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5367 _17044_/Q vssd1 vssd1 vccd1 vccd1 hold5367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4633 _17646_/Q vssd1 vssd1 vccd1 vccd1 hold4633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5378 _09934_/X vssd1 vssd1 vccd1 vccd1 _16468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4644 _12214_/X vssd1 vssd1 vccd1 vccd1 _17228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5389 _16889_/Q vssd1 vssd1 vccd1 vccd1 hold5389/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3910 hold5844/X vssd1 vssd1 vccd1 vccd1 hold5845/A sky130_fd_sc_hd__buf_4
Xhold4655 _17225_/Q vssd1 vssd1 vccd1 vccd1 hold4655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4666 _10429_/X vssd1 vssd1 vccd1 vccd1 _16633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3921 _13852_/Y vssd1 vssd1 vccd1 vccd1 _17737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3932 _13878_/Y vssd1 vssd1 vccd1 vccd1 _13879_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4677 _17265_/Q vssd1 vssd1 vccd1 vccd1 hold4677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3943 _12336_/Y vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4688 _16418_/Q vssd1 vssd1 vccd1 vccd1 hold4688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3954 _11797_/Y vssd1 vssd1 vccd1 vccd1 _17089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4699 _10180_/X vssd1 vssd1 vccd1 vccd1 _16550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3965 _16594_/Q vssd1 vssd1 vccd1 vccd1 hold3965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3976 _16571_/Q vssd1 vssd1 vccd1 vccd1 hold3976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3987 _16753_/Q vssd1 vssd1 vccd1 vccd1 hold3987/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout155 _13001_/S vssd1 vssd1 vccd1 vccd1 _12953_/S sky130_fd_sc_hd__clkbuf_8
Xfanout166 _13823_/B vssd1 vssd1 vccd1 vccd1 _13862_/B sky130_fd_sc_hd__buf_2
Xhold3998 _13342_/X vssd1 vssd1 vccd1 vccd1 _17567_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout177 _11741_/B vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__buf_4
Xfanout188 _12362_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__buf_4
Xfanout199 fanout209/X vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__clkbuf_4
X_07989_ hold2707/X _07991_/A2 _07988_/X _08143_/A vssd1 vssd1 vccd1 vccd1 _07989_/X
+ sky130_fd_sc_hd__o211a_1
X_09728_ _18313_/Q hold5635/X _11201_/C vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__mux2_1
X_09659_ hold775/X hold3386/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__mux2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12670_ hold1857/X _17401_/Q _12679_/S vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18204_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ hold2038/X hold4860/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18373_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ hold300/A hold273/A vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__or2_1
XFILLER_0_53_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11552_ _17856_/Q hold4469/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10503_ _10521_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__or2_1
X_11483_ hold1288/X _16985_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__mux2_1
X_14271_ hold886/X _14272_/B _14270_/Y _14388_/A vssd1 vssd1 vccd1 vccd1 hold887/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _18417_/CLK _16010_/D vssd1 vssd1 vccd1 vccd1 _16010_/Q sky130_fd_sc_hd__dfxtp_1
X_10434_ _10485_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13222_ _13222_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13153_ _13153_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__and2_1
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ _11097_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ hold1375/X hold4739/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__mux2_1
X_17961_ _18055_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
X_13084_ hold3610/X _13083_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_1
Xhold5890 _18459_/Q vssd1 vssd1 vccd1 vccd1 hold5890/X sky130_fd_sc_hd__dlygate4sd3_1
X_10296_ _10551_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10296_/X sky130_fd_sc_hd__or2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12035_ hold2222/X hold4704/X _12329_/C vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__mux2_1
X_16912_ _17856_/CLK _16912_/D vssd1 vssd1 vccd1 vccd1 _16912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17892_ _17892_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_1
X_16843_ _18046_/CLK _16843_/D vssd1 vssd1 vccd1 vccd1 _16843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ _18009_/CLK _16774_/D vssd1 vssd1 vccd1 vccd1 _16774_/Q sky130_fd_sc_hd__dfxtp_1
X_13986_ _14774_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_279_wb_clk_i clkbuf_5_18__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17923_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15725_ _17731_/CLK hold923/X vssd1 vssd1 vccd1 vccd1 hold922/A sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12937_ hold1416/X _17490_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_208_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17898_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _18456_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
X_15656_ _17232_/CLK _15656_/D vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ hold1073/X hold3281/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__mux2_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ hold939/X _14612_/B _14606_/Y _14807_/C1 vssd1 vssd1 vccd1 vccd1 hold940/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18375_ _18416_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
X_11819_ hold2550/X hold3811/X _12299_/C vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__mux2_1
X_15587_ _17865_/CLK _15587_/D vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ hold1950/X _17444_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ _18425_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _17326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14538_ hold2012/X _14541_/B _14537_/Y _13913_/A vssd1 vssd1 vccd1 vccd1 _14538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17257_ _17257_/CLK _17257_/D vssd1 vssd1 vccd1 vccd1 _17257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14469_ hold747/X _14479_/B vssd1 vssd1 vccd1 vccd1 _14469_/X sky130_fd_sc_hd__or2_1
X_16208_ _17439_/CLK _16208_/D vssd1 vssd1 vccd1 vccd1 _16208_/Q sky130_fd_sc_hd__dfxtp_1
X_17188_ _17844_/CLK _17188_/D vssd1 vssd1 vccd1 vccd1 _17188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _17314_/CLK _16139_/D vssd1 vssd1 vccd1 vccd1 hold659/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3206 _16579_/Q vssd1 vssd1 vccd1 vccd1 hold3206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3217 _17592_/Q vssd1 vssd1 vccd1 vccd1 hold3217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ hold59/X _16098_/Q _08997_/S vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__mux2_1
Xhold3228 _17482_/Q vssd1 vssd1 vccd1 vccd1 hold3228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3239 _10519_/X vssd1 vssd1 vccd1 vccd1 _16663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2505 _17812_/Q vssd1 vssd1 vccd1 vccd1 hold2505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 _15618_/Q vssd1 vssd1 vccd1 vccd1 hold2516/X sky130_fd_sc_hd__dlygate4sd3_1
X_07912_ _14529_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07912_/X sky130_fd_sc_hd__or2_1
Xhold2527 _08414_/X vssd1 vssd1 vccd1 vccd1 _15837_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08892_ hold136/X hold555/X _08930_/S vssd1 vssd1 vccd1 vccd1 hold556/A sky130_fd_sc_hd__mux2_1
Xhold2538 _18031_/Q vssd1 vssd1 vccd1 vccd1 hold2538/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 _18077_/Q vssd1 vssd1 vccd1 vccd1 hold1804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 _15528_/X vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 _14571_/X vssd1 vssd1 vccd1 vccd1 _18080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 _15633_/Q vssd1 vssd1 vccd1 vccd1 hold1826/X sky130_fd_sc_hd__dlygate4sd3_1
X_07843_ _15521_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07843_/X sky130_fd_sc_hd__or2_1
Xhold1837 _14727_/X vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1848 _15713_/Q vssd1 vssd1 vccd1 vccd1 hold1848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _15746_/Q vssd1 vssd1 vccd1 vccd1 hold1859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09513_ _11067_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09444_ _09447_/B _09447_/C _09447_/D vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__and3_1
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _15471_/A _09375_/B _09375_/C _09375_/D vssd1 vssd1 vccd1 vccd1 _09375_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08326_ hold1934/X _08323_/B _08325_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08326_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ hold1650/X _08262_/B _08256_/X _08257_/C1 vssd1 vssd1 vccd1 vccd1 _08257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ hold2854/X _08209_/B _08187_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _08188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5120 _16378_/Q vssd1 vssd1 vccd1 vccd1 hold5120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5131 _13363_/X vssd1 vssd1 vccd1 vccd1 _17574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5142 _16676_/Q vssd1 vssd1 vccd1 vccd1 hold5142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5153 _09979_/X vssd1 vssd1 vccd1 vccd1 _16483_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5164 _17610_/Q vssd1 vssd1 vccd1 vccd1 hold5164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5175 _16449_/Q vssd1 vssd1 vccd1 vccd1 hold5175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4430 _11461_/X vssd1 vssd1 vccd1 vccd1 _16977_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10150_ hold3349/X _10646_/B _10149_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10150_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5186 _15353_/X vssd1 vssd1 vccd1 vccd1 _15354_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4441 _16976_/Q vssd1 vssd1 vccd1 vccd1 hold4441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4452 _10954_/X vssd1 vssd1 vccd1 vccd1 _16808_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5197 _16645_/Q vssd1 vssd1 vccd1 vccd1 hold5197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4463 _17666_/Q vssd1 vssd1 vccd1 vccd1 hold4463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4474 _10933_/X vssd1 vssd1 vccd1 vccd1 _16801_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4485 _09886_/X vssd1 vssd1 vccd1 vccd1 _16452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3740 _17122_/Q vssd1 vssd1 vccd1 vccd1 hold3740/X sky130_fd_sc_hd__dlygate4sd3_1
X_10081_ hold4777/X _10571_/B _10080_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _10081_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4496 _17597_/Q vssd1 vssd1 vccd1 vccd1 hold4496/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3751 _16712_/Q vssd1 vssd1 vccd1 vccd1 hold3751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3762 _16399_/Q vssd1 vssd1 vccd1 vccd1 hold3762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3773 _17102_/Q vssd1 vssd1 vccd1 vccd1 hold3773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3784 _16726_/Q vssd1 vssd1 vccd1 vccd1 hold3784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3795 _13843_/Y vssd1 vssd1 vccd1 vccd1 _17734_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13840_ _13873_/A _13840_/B vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13771_ hold4471/X _13868_/B _13770_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13771_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_301_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17726_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10983_ _11658_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__or2_1
X_15510_ hold5977/X _15560_/A2 hold945/X _12885_/A vssd1 vssd1 vccd1 vccd1 hold946/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ hold3512/X _12721_/X _12806_/S vssd1 vssd1 vccd1 vccd1 _12723_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _18243_/CLK _16490_/D vssd1 vssd1 vccd1 vccd1 _16490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15441_ hold398/X _09392_/D _09386_/D hold339/X _15436_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/D sky130_fd_sc_hd__a221o_1
X_12653_ hold3102/X _12652_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18160_ _18232_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
X_11604_ _12153_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15372_ _15489_/A _15372_/B _15372_/C _15372_/D vssd1 vssd1 vccd1 vccd1 _15372_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12584_ hold2925/X _12583_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17111_ _17779_/CLK _17111_/D vssd1 vssd1 vccd1 vccd1 _17111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14323_ hold2304/X _14326_/B _14322_/Y _14384_/A vssd1 vssd1 vccd1 vccd1 _14323_/X
+ sky130_fd_sc_hd__o211a_1
X_18091_ _18219_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
X_11535_ _11631_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__or2_1
XFILLER_0_108_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17042_ _17890_/CLK _17042_/D vssd1 vssd1 vccd1 vccd1 _17042_/Q sky130_fd_sc_hd__dfxtp_1
X_14254_ _14988_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11658_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13205_ _13204_/X hold3135/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__mux2_1
X_10417_ hold4057/X _10631_/B _10416_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10417_/X
+ sky130_fd_sc_hd__o211a_1
X_11397_ _12036_/A _11397_/B vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__or2_1
X_14185_ hold804/X _14202_/B _14184_/X _14548_/C1 vssd1 vssd1 vccd1 vccd1 hold805/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13136_ _13129_/X _13135_/X _13312_/B1 vssd1 vssd1 vccd1 vccd1 _17535_/D sky130_fd_sc_hd__o21a_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10348_ hold4254/X _11213_/B _10347_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ hold4883/X _10568_/B _10278_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _10279_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13066_/X _16901_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__mux2_1
X_17944_ _18043_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12018_ _12018_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__or2_1
X_17875_ _17904_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _18066_/CLK _16826_/D vssd1 vssd1 vccd1 vccd1 _16826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16757_ _18158_/CLK _16757_/D vssd1 vssd1 vccd1 vccd1 _16757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13969_ hold1889/X _13980_/B _13968_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _13969_/X
+ sky130_fd_sc_hd__o211a_1
X_15708_ _17276_/CLK _15708_/D vssd1 vssd1 vccd1 vccd1 hold369/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16688_ _18118_/CLK _16688_/D vssd1 vssd1 vccd1 vccd1 _16688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _17282_/CLK _15639_/D vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18427_ _18427_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _15543_/A _09164_/B vssd1 vssd1 vccd1 vccd1 _09160_/Y sky130_fd_sc_hd__nand2_1
X_18358_ _18358_/CLK hold807/X vssd1 vssd1 vccd1 vccd1 hold806/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__and2_1
X_17309_ _17329_/CLK _17309_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ hold1482/X _09106_/B _09090_/X _14364_/A vssd1 vssd1 vccd1 vccd1 _09091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18289_ _18353_/CLK hold836/X vssd1 vssd1 vccd1 vccd1 hold835/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ hold2441/X _08033_/B _08041_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _08042_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold901 hold901/A vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__clkbuf_2
Xhold912 hold912/A vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/A vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold934 hold934/A vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 hold945/A vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 hold967/A vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__buf_4
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3003 _16230_/Q vssd1 vssd1 vccd1 vccd1 hold3003/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3014 _17388_/Q vssd1 vssd1 vccd1 vccd1 hold3014/X sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _13094_/A _10779_/A _09992_/X vssd1 vssd1 vccd1 vccd1 _09993_/Y sky130_fd_sc_hd__a21oi_1
Xhold3025 _17427_/Q vssd1 vssd1 vccd1 vccd1 hold3025/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3036 _12743_/X vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2302 _17372_/Q vssd1 vssd1 vccd1 vccd1 hold2302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3047 _12521_/X vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08944_ _12402_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _16089_/D sky130_fd_sc_hd__and2_1
Xhold2313 _14542_/X vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3058 _12971_/X vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 _17408_/Q vssd1 vssd1 vccd1 vccd1 hold3069/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 _18006_/Q vssd1 vssd1 vccd1 vccd1 hold2324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2335 _07832_/X vssd1 vssd1 vccd1 vccd1 _15561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2346 _18397_/Q vssd1 vssd1 vccd1 vccd1 hold2346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1601 hold6014/X vssd1 vssd1 vccd1 vccd1 hold1601/X sky130_fd_sc_hd__buf_1
Xhold1612 _18215_/Q vssd1 vssd1 vccd1 vccd1 hold1612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 _18449_/Q vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08875_ _15334_/A hold455/X vssd1 vssd1 vccd1 vccd1 _16055_/D sky130_fd_sc_hd__and2_1
Xhold1623 hold6036/X vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__buf_1
Xhold2368 _15538_/X vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 _18175_/Q vssd1 vssd1 vccd1 vccd1 hold2379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 _15727_/Q vssd1 vssd1 vccd1 vccd1 hold1634/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1645 _08457_/X vssd1 vssd1 vccd1 vccd1 _15857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07826_ _07826_/A _13048_/A vssd1 vssd1 vccd1 vccd1 _07826_/X sky130_fd_sc_hd__and2_1
Xhold1656 _18300_/Q vssd1 vssd1 vccd1 vccd1 hold1656/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1667 _16152_/Q vssd1 vssd1 vccd1 vccd1 hold1667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 _08057_/X vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1689 _14833_/X vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _07785_/Y _09472_/B _15314_/A _09426_/X vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09358_ _09400_/A _09363_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09358_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_63_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08309_ _15533_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08309_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09289_ _14970_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09289_/X sky130_fd_sc_hd__or2_1
X_11320_ hold5003/X _11798_/B _11319_/X _13941_/A vssd1 vssd1 vccd1 vccd1 _11320_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11251_ hold4540/X _11732_/B _11250_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ hold2277/X hold4891/X _10628_/C vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__mux2_1
X_11182_ _11194_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__nor2_1
Xhold4260 _13546_/X vssd1 vssd1 vccd1 vccd1 _17635_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10133_ hold1809/X _16535_/Q _10523_/S vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__mux2_1
Xhold4271 _16622_/Q vssd1 vssd1 vccd1 vccd1 hold4271/X sky130_fd_sc_hd__dlygate4sd3_1
X_15990_ _17524_/CLK _15990_/D vssd1 vssd1 vccd1 vccd1 hold694/A sky130_fd_sc_hd__dfxtp_1
Xhold4282 _13348_/X vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4293 _16389_/Q vssd1 vssd1 vccd1 vccd1 hold4293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3570 _17704_/Q vssd1 vssd1 vccd1 vccd1 hold3570/X sky130_fd_sc_hd__dlygate4sd3_1
X_10064_ _16512_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__and3_1
Xhold3581 _17357_/Q vssd1 vssd1 vccd1 vccd1 hold3581/X sky130_fd_sc_hd__dlygate4sd3_1
X_14941_ hold1671/X _14952_/B _14940_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14941_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3592 _17487_/Q vssd1 vssd1 vccd1 vccd1 hold3592/X sky130_fd_sc_hd__dlygate4sd3_1
X_17660_ _17723_/CLK _17660_/D vssd1 vssd1 vccd1 vccd1 _17660_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2880 _18118_/Q vssd1 vssd1 vccd1 vccd1 hold2880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2891 _18223_/Q vssd1 vssd1 vccd1 vccd1 hold2891/X sky130_fd_sc_hd__dlygate4sd3_1
X_14872_ hold735/X _14894_/B vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__or2_1
X_16611_ _18230_/CLK _16611_/D vssd1 vssd1 vccd1 vccd1 _16611_/Q sky130_fd_sc_hd__dfxtp_1
X_13823_ _17728_/Q _13823_/B _13862_/C vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__and3_1
X_17591_ _17719_/CLK _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16542_ _18222_/CLK _16542_/D vssd1 vssd1 vccd1 vccd1 _16542_/Q sky130_fd_sc_hd__dfxtp_1
X_13754_ hold1891/X _17705_/Q _13880_/C vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__mux2_1
X_10966_ hold5576/X _11156_/B _10965_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12705_ _12777_/A _12705_/B vssd1 vssd1 vccd1 vccd1 _17411_/D sky130_fd_sc_hd__and2_1
X_16473_ _18358_/CLK _16473_/D vssd1 vssd1 vccd1 vccd1 _16473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13685_ hold1650/X hold5092/X _13880_/C vssd1 vssd1 vccd1 vccd1 _13686_/B sky130_fd_sc_hd__mux2_1
X_10897_ hold3915/X _10897_/A2 _10896_/X _14733_/C1 vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__o211a_1
X_18212_ _18266_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
X_15424_ _15473_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__and2_1
XFILLER_0_183_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ _12855_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _17388_/D sky130_fd_sc_hd__and2_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18143_ _18267_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
X_15355_ _15355_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12567_ _12996_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _17365_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ _14986_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__or2_1
X_11518_ hold4767/X _11741_/B _11517_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11518_/X
+ sky130_fd_sc_hd__o211a_1
X_18074_ _18080_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
X_15286_ _17332_/Q _15486_/B1 _15485_/B1 hold354/X vssd1 vssd1 vccd1 vccd1 _15286_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12498_ _17342_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__or2_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 hold546/X vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__buf_4
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17025_ _17873_/CLK _17025_/D vssd1 vssd1 vccd1 vccd1 _17025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ hold1517/X _14266_/B _14236_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14237_/X
+ sky130_fd_sc_hd__o211a_1
X_11449_ hold4178/X _11735_/B _11448_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14168_ _14740_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14168_/X sky130_fd_sc_hd__or2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13119_ _13183_/A1 _13117_/X _13118_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13119_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_294_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14099_ hold1353/X _14105_/A2 _14098_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14099_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _18236_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_223_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17779_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08660_ _12426_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _15952_/D sky130_fd_sc_hd__and2_1
X_17858_ _17889_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
X_16809_ _18047_/CLK _16809_/D vssd1 vssd1 vccd1 vccd1 _16809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ _15344_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__and2_1
X_17789_ _18051_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _15541_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ hold2457/X _09177_/A2 _09142_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _09143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ _15515_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08025_ _15539_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout2 fanout2/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_4
XFILLER_0_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 hold720/A vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 hold731/A vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 hold764/A vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold775 hold775/A vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold877/X vssd1 vssd1 vccd1 vccd1 hold878/A sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ hold4913/X _10070_/B _09975_/X _15028_/A vssd1 vssd1 vccd1 vccd1 _09976_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2110 _07870_/X vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2121 _16201_/Q vssd1 vssd1 vccd1 vccd1 hold2121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2132 _08208_/X vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08927_ _12438_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _16081_/D sky130_fd_sc_hd__and2_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2143 _15689_/Q vssd1 vssd1 vccd1 vccd1 hold2143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2154 _08485_/X vssd1 vssd1 vccd1 vccd1 _15871_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _16272_/Q vssd1 vssd1 vccd1 vccd1 hold2165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1420 _17515_/Q vssd1 vssd1 vccd1 vccd1 hold1420/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1431 _14947_/X vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2176 _12512_/X vssd1 vssd1 vccd1 vccd1 hold2176/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1442 _15694_/Q vssd1 vssd1 vccd1 vccd1 hold1442/X sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ hold44/X hold321/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__mux2_1
Xhold2187 _18117_/Q vssd1 vssd1 vccd1 vccd1 hold2187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1453 _15535_/A vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2198 _14039_/X vssd1 vssd1 vccd1 vccd1 _17825_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 _14265_/X vssd1 vssd1 vccd1 vccd1 _17933_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1475 _17939_/Q vssd1 vssd1 vccd1 vccd1 hold1475/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1486 _18331_/Q vssd1 vssd1 vccd1 vccd1 hold1486/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _18459_/Q _18460_/Q vssd1 vssd1 vccd1 vccd1 _07809_/X sky130_fd_sc_hd__or2_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _15669_/Q vssd1 vssd1 vccd1 vccd1 hold1497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ hold380/X _16015_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold381/A sky130_fd_sc_hd__mux2_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ hold2427/X _16764_/Q _11210_/C vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__mux2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ hold1197/X hold5423/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13470_ _13779_/A _13470_/B vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ hold2936/X hold5312/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10683_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ hold5/X hold398/X _12443_/S vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15140_ hold2981/X hold609/X _15139_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15140_/X
+ sky130_fd_sc_hd__o211a_1
X_12352_ _13888_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ hold402/X hold3613/X _12329_/C vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__mux2_1
X_15071_ _15233_/A hold2196/X hold302/X vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__mux2_1
X_12283_ hold4635/X _12377_/B _12282_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _12283_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _15529_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__or2_1
X_11234_ hold1780/X hold4852/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__mux2_1
X_11165_ _16879_/Q _11171_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__and3_1
XFILLER_0_140_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4090 _13702_/X vssd1 vssd1 vccd1 vccd1 _17687_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10116_ _10524_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__or2_1
X_15973_ _17292_/CLK _15973_/D vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
X_11096_ hold2848/X _16856_/Q _11192_/C vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _13238_/A _09975_/A _10046_/X vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__a21oi_1
X_17712_ _17743_/CLK _17712_/D vssd1 vssd1 vccd1 vccd1 _17712_/Q sky130_fd_sc_hd__dfxtp_1
X_14924_ _15193_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__or2_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold4/X vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
X_17643_ _17734_/CLK _17643_/D vssd1 vssd1 vccd1 vccd1 _17643_/Q sky130_fd_sc_hd__dfxtp_1
X_14855_ hold2507/X _14882_/B _14854_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14855_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ hold3865/X _13710_/A _13805_/X vssd1 vssd1 vccd1 vccd1 _13806_/Y sky130_fd_sc_hd__a21oi_1
X_17574_ _17736_/CLK _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14786_ _14786_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14786_/X sky130_fd_sc_hd__or2_1
X_11998_ hold4797/X _12320_/B _11997_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16525_ _18266_/CLK _16525_/D vssd1 vssd1 vccd1 vccd1 _16525_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _13737_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__or2_1
XFILLER_0_156_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10949_ hold2338/X _16807_/Q _11156_/C vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ _18273_/CLK _16456_/D vssd1 vssd1 vccd1 vccd1 _16456_/Q sky130_fd_sc_hd__dfxtp_1
X_13668_ _13764_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _17316_/Q _09357_/A _15484_/B1 hold373/X _15406_/X vssd1 vssd1 vccd1 vccd1
+ _15412_/B sky130_fd_sc_hd__a221o_1
X_12619_ hold2934/X _17384_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__mux2_1
X_16387_ _18388_/CLK _16387_/D vssd1 vssd1 vccd1 vccd1 _16387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13599_ _13779_/A _13599_/B vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18126_ _18126_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_1
X_15338_ hold168/X _15484_/A2 _15451_/A2 hold186/X vssd1 vssd1 vccd1 vccd1 _15338_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5708 _11476_/X vssd1 vssd1 vccd1 vccd1 _16982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5719 _16815_/Q vssd1 vssd1 vccd1 vccd1 hold5719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _18061_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
X_15269_ hold559/X _09365_/B _09392_/C hold538/X _15268_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17008_ _17856_/CLK _17008_/D vssd1 vssd1 vccd1 vccd1 _17008_/Q sky130_fd_sc_hd__dfxtp_1
X_09830_ hold2381/X hold3307/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__mux2_1
Xfanout507 _10610_/C vssd1 vssd1 vccd1 vccd1 _10646_/C sky130_fd_sc_hd__clkbuf_8
Xfanout518 _10649_/C vssd1 vssd1 vccd1 vccd1 _10640_/C sky130_fd_sc_hd__clkbuf_8
Xfanout529 _09277_/S vssd1 vssd1 vccd1 vccd1 _09283_/S sky130_fd_sc_hd__clkbuf_8
X_09761_ hold1523/X hold5009/X _10055_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__mux2_1
X_08712_ _15473_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _15977_/D sky130_fd_sc_hd__and2_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ hold3060/X _16388_/Q _10022_/C vssd1 vssd1 vccd1 vccd1 _09693_/B sky130_fd_sc_hd__mux2_1
X_08643_ hold140/X hold712/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ hold8/X hold164/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__mux2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ _14218_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ _15344_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _16145_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ hold2449/X _08029_/B _08007_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _08008_/X
+ sky130_fd_sc_hd__o211a_1
Xhold550 hold550/A vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_145_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold572 input50/X vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold583 input56/X vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 hold594/A vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ hold1004/X _16477_/Q _10601_/C vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__mux2_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ hold1465/X _17501_/Q _12982_/S vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__mux2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 _14133_/X vssd1 vssd1 vccd1 vccd1 _17870_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 input40/X vssd1 vssd1 vccd1 vccd1 hold1261/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ hold2805/X hold5028/X _12305_/C vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__mux2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _08328_/X vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _08198_/X vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _18003_/Q vssd1 vssd1 vccd1 vccd1 hold1294/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14980_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__or2_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ hold2630/X hold3174/X _12332_/C vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__mux2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _11097_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__or2_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14980_/A _14557_/Y hold1814/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _14571_/X
+ sky130_fd_sc_hd__o211a_1
X_11783_ _17085_/Q _11783_/B _11783_/C vssd1 vssd1 vccd1 vccd1 _11783_/X sky130_fd_sc_hd__and3_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16310_ _17511_/CLK _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/Q sky130_fd_sc_hd__dfxtp_1
X_13522_ hold4787/X _13805_/B _13521_/X _12756_/A vssd1 vssd1 vccd1 vccd1 _13522_/X
+ sky130_fd_sc_hd__o211a_1
X_17290_ _17313_/CLK _17290_/D vssd1 vssd1 vccd1 vccd1 hold578/A sky130_fd_sc_hd__dfxtp_1
X_10734_ _11103_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ _17428_/CLK _16241_/D vssd1 vssd1 vccd1 vccd1 _16241_/Q sky130_fd_sc_hd__dfxtp_1
X_13453_ hold4651/X _13856_/B _13452_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ _11637_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _15354_/A hold562/X vssd1 vssd1 vccd1 vccd1 _17295_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16172_ _17517_/CLK _16172_/D vssd1 vssd1 vccd1 vccd1 _16172_/Q sky130_fd_sc_hd__dfxtp_1
X_13384_ hold4377/X _13823_/B _13383_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _13384_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10596_ _16529_/Q _10524_/A _10595_/X vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ _15123_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__or2_1
X_12335_ _17269_/Q _12341_/B _12341_/C vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15054_ _15054_/A hold266/X vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ hold1966/X hold4718/X _12356_/C vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ hold1035/X _14036_/B _14004_/X _13939_/A vssd1 vssd1 vccd1 vccd1 _14005_/X
+ sky130_fd_sc_hd__o211a_1
X_11217_ hold5248/X _11121_/A _11216_/X vssd1 vssd1 vccd1 vccd1 _11217_/Y sky130_fd_sc_hd__a21oi_1
X_12197_ hold1920/X _17223_/Q _12308_/C vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput81 _13201_/A vssd1 vssd1 vccd1 vccd1 output81/X sky130_fd_sc_hd__buf_6
Xoutput92 _13281_/A vssd1 vssd1 vccd1 vccd1 output92/X sky130_fd_sc_hd__buf_6
X_11148_ hold3607/X _11061_/A _11147_/X vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__a21oi_1
X_15956_ _17302_/CLK _15956_/D vssd1 vssd1 vccd1 vccd1 hold416/A sky130_fd_sc_hd__dfxtp_1
X_11079_ _11658_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__or2_1
X_14907_ hold5952/X hold657/A _14906_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 hold658/A
+ sky130_fd_sc_hd__o211a_1
X_15887_ _18425_/CLK _15887_/D vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17626_ _17725_/CLK _17626_/D vssd1 vssd1 vccd1 vccd1 _17626_/Q sky130_fd_sc_hd__dfxtp_1
X_14838_ _15123_/A _14838_/B vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__or2_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ _18229_/CLK _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
X_14769_ hold2379/X _14774_/B _14768_/Y _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14769_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16508_ _18389_/CLK _16508_/D vssd1 vssd1 vccd1 vccd1 _16508_/Q sky130_fd_sc_hd__dfxtp_1
X_08290_ hold2997/X _08323_/B _08289_/X _08351_/A vssd1 vssd1 vccd1 vccd1 _08290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17488_ _17516_/CLK _17488_/D vssd1 vssd1 vccd1 vccd1 _17488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16439_ _18388_/CLK _16439_/D vssd1 vssd1 vccd1 vccd1 _16439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5505 _11560_/X vssd1 vssd1 vccd1 vccd1 _17010_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18109_ _18267_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5516 _16393_/Q vssd1 vssd1 vccd1 vccd1 hold5516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5527 _10930_/X vssd1 vssd1 vccd1 vccd1 _16800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5538 _16863_/Q vssd1 vssd1 vccd1 vccd1 hold5538/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4804 _11938_/X vssd1 vssd1 vccd1 vccd1 _17136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5549 _10867_/X vssd1 vssd1 vccd1 vccd1 _16779_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4815 _16900_/Q vssd1 vssd1 vccd1 vccd1 hold4815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4826 _17638_/Q vssd1 vssd1 vccd1 vccd1 hold4826/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4837 _13420_/X vssd1 vssd1 vccd1 vccd1 _17593_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4848 _17711_/Q vssd1 vssd1 vccd1 vccd1 hold4848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4859 _10177_/X vssd1 vssd1 vccd1 vccd1 _16549_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout304 _09981_/A vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__buf_2
Xfanout315 _10560_/A vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__buf_4
Xfanout326 _09951_/A vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__buf_4
Xfanout337 _09493_/Y vssd1 vssd1 vccd1 vccd1 fanout337/X sky130_fd_sc_hd__buf_8
X_09813_ _09933_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__or2_1
Xfanout348 _08997_/S vssd1 vssd1 vccd1 vccd1 _08993_/S sky130_fd_sc_hd__buf_8
Xfanout359 _08562_/S vssd1 vssd1 vccd1 vccd1 _08590_/S sky130_fd_sc_hd__buf_8
XFILLER_0_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _09933_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _11082_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _09011_/A _08626_/B vssd1 vssd1 vccd1 vccd1 _15935_/D sky130_fd_sc_hd__and2_1
XFILLER_0_179_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _15284_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _15902_/D sky130_fd_sc_hd__and2_1
XFILLER_0_167_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08488_ _14774_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ hold4361/X _10640_/B _10449_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ hold2544/X _09106_/B _09108_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _09109_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ hold3502/X _10571_/B _10380_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _10381_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _13794_/A _12120_/B vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _12051_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__or2_1
Xhold380 hold62/X vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__buf_4
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold391 hold391/A vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ hold5584/X _11213_/B _11001_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _11002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout860 hold1550/X vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__buf_4
Xfanout871 _15221_/A vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__clkbuf_16
X_15810_ _17428_/CLK _15810_/D vssd1 vssd1 vccd1 vccd1 _15810_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout882 hold967/X vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__buf_4
X_16790_ _18025_/CLK _16790_/D vssd1 vssd1 vccd1 vccd1 _16790_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout893 hold490/X vssd1 vssd1 vccd1 vccd1 _14511_/A sky130_fd_sc_hd__buf_8
X_15741_ _17743_/CLK _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ hold3583/X _12952_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12954_/B sky130_fd_sc_hd__mux2_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 _14059_/X vssd1 vssd1 vccd1 vccd1 _17834_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 _18337_/Q vssd1 vssd1 vccd1 vccd1 hold1091/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11904_ _13797_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _17253_/CLK hold968/X vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18046_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18460_ _18460_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ hold3023/X _12883_/X _12911_/S vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__mux2_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ hold1811/X _14610_/B _14622_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _14623_/X
+ sky130_fd_sc_hd__o211a_1
X_17411_ _17435_/CLK _17411_/D vssd1 vssd1 vccd1 vccd1 _17411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _12267_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__or2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _18391_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17342_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _17342_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ hold5966/X _14554_/A2 _14553_/X _14352_/A vssd1 vssd1 vccd1 vccd1 hold852/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ hold5331/X _11670_/A _11765_/X vssd1 vssd1 vccd1 vccd1 _11766_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ hold2383/X _17622_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__mux2_1
X_17273_ _17583_/CLK _17273_/D vssd1 vssd1 vccd1 vccd1 _17273_/Q sky130_fd_sc_hd__dfxtp_1
X_10717_ hold5450/X _11762_/B _10716_/X _13913_/A vssd1 vssd1 vccd1 vccd1 _10717_/X
+ sky130_fd_sc_hd__o211a_1
X_14485_ _15545_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11697_ _11697_/A _11697_/B vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16224_ _17456_/CLK _16224_/D vssd1 vssd1 vccd1 vccd1 _16224_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ hold2562/X hold3997/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13437_/B sky130_fd_sc_hd__mux2_1
X_10648_ _11218_/A _10648_/B vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_181_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16155_ _17494_/CLK _16155_/D vssd1 vssd1 vccd1 vccd1 _16155_/Q sky130_fd_sc_hd__dfxtp_1
X_13367_ hold1397/X hold3196/X _13388_/S vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__mux2_1
X_10579_ _10588_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15106_ hold1091/X _15109_/B _15105_/X _15172_/C1 vssd1 vssd1 vccd1 vccd1 _15106_/X
+ sky130_fd_sc_hd__o211a_1
X_12318_ hold3825/X _12267_/A _12317_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__a21oi_1
X_16086_ _17329_/CLK _16086_/D vssd1 vssd1 vccd1 vccd1 hold396/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ _17588_/Q _17122_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _14984_/A hold2771/X hold302/X vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_139_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ _13749_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2709 _17994_/Q vssd1 vssd1 vccd1 vccd1 hold2709/X sky130_fd_sc_hd__dlygate4sd3_1
X_07790_ hold270/X vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__inv_2
X_16988_ _17900_/CLK _16988_/D vssd1 vssd1 vccd1 vccd1 _16988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15939_ _18417_/CLK _15939_/D vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09460_ _09463_/C _09463_/D _09463_/B vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_176_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ _15525_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08411_/X sky130_fd_sc_hd__or2_1
X_17609_ _17649_/CLK _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_1
X_09391_ hold5853/A _09342_/B _09342_/Y _09390_/X _12442_/A vssd1 vssd1 vccd1 vccd1
+ _09391_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08342_ hold756/X hold910/X _08390_/S vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ hold1509/X _08268_/B _08272_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _08273_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6003 data_in[28] vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6014 _16323_/Q vssd1 vssd1 vccd1 vccd1 hold6014/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6025 data_in[1] vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6036 _16314_/Q vssd1 vssd1 vccd1 vccd1 hold6036/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5302 _11227_/Y vssd1 vssd1 vccd1 vccd1 _16899_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5313 _11163_/Y vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5324 _16918_/Q vssd1 vssd1 vccd1 vccd1 hold5324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5335 _11497_/X vssd1 vssd1 vccd1 vccd1 _16989_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4601 _17052_/Q vssd1 vssd1 vccd1 vccd1 hold4601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5346 _16823_/Q vssd1 vssd1 vccd1 vccd1 hold5346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5357 _11769_/Y vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4612 _11347_/X vssd1 vssd1 vccd1 vccd1 _16939_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4623 _17193_/Q vssd1 vssd1 vccd1 vccd1 hold4623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5368 _11566_/X vssd1 vssd1 vccd1 vccd1 _17012_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5379 _16433_/Q vssd1 vssd1 vccd1 vccd1 hold5379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4634 _13483_/X vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3900 _16346_/Q vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__buf_1
XFILLER_0_160_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4645 _16884_/Q vssd1 vssd1 vccd1 vccd1 hold4645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3911 _09385_/X vssd1 vssd1 vccd1 vccd1 _16281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4656 _12109_/X vssd1 vssd1 vccd1 vccd1 _17193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4667 _17280_/Q vssd1 vssd1 vccd1 vccd1 hold4667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3922 _16796_/Q vssd1 vssd1 vccd1 vccd1 hold3922/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3933 _13879_/Y vssd1 vssd1 vccd1 vccd1 _17746_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4678 _12229_/X vssd1 vssd1 vccd1 vccd1 _17233_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4689 _09688_/X vssd1 vssd1 vccd1 vccd1 _16386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3944 _12337_/Y vssd1 vssd1 vccd1 vccd1 _17269_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3955 _16002_/Q vssd1 vssd1 vccd1 vccd1 _15325_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3966 _10216_/X vssd1 vssd1 vccd1 vccd1 _16562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3977 _10147_/X vssd1 vssd1 vccd1 vccd1 _16539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout156 _12980_/S vssd1 vssd1 vccd1 vccd1 _13001_/S sky130_fd_sc_hd__buf_6
Xfanout167 _13823_/B vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__buf_4
Xhold3988 _10693_/X vssd1 vssd1 vccd1 vccd1 _16721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3999 _16395_/Q vssd1 vssd1 vccd1 vccd1 hold3999/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout178 _11741_/B vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__buf_4
X_07988_ _15557_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
Xfanout189 _12362_/B vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__buf_4
X_09727_ hold5433/X _10013_/B _09726_/X _15058_/A vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__o211a_1
X_09658_ hold4357/X _11177_/B _09657_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _09658_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ hold41/X hold551/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ hold3484/X _10067_/B _09588_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09589_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ hold5096/X _12305_/B _11619_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11620_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11551_ hold4663/X _12323_/B _11550_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ hold2507/X hold3972/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__mux2_1
X_14270_ _14950_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__nand2_1
X_11482_ hold4579/X _11798_/B _11481_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _11482_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_160_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18198_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13220_/X hold3619/X _13309_/S vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__mux2_1
X_10433_ hold2774/X hold4061/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_104_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _13145_/X _13151_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17537_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10364_ hold2746/X _16612_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__mux2_1
X_12103_ hold4443/X _12302_/B _12102_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _12103_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5880 hold6001/X vssd1 vssd1 vccd1 vccd1 _18463_/A sky130_fd_sc_hd__clkbuf_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13082_/X _16903_/Q _13251_/S vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux2_1
X_17960_ _18158_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
X_10295_ hold2363/X hold3334/X _10589_/C vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__mux2_1
Xhold5891 _07793_/X vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__dlygate4sd3_1
X_12034_ hold4985/X _12311_/B _12033_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _12034_/X
+ sky130_fd_sc_hd__o211a_1
X_16911_ _17887_/CLK _16911_/D vssd1 vssd1 vccd1 vccd1 _16911_/Q sky130_fd_sc_hd__dfxtp_1
X_17891_ _17891_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_1
X_16842_ _18013_/CLK _16842_/D vssd1 vssd1 vccd1 vccd1 _16842_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout690 _12951_/A vssd1 vssd1 vccd1 vccd1 _12996_/A sky130_fd_sc_hd__buf_4
X_13985_ hold2125/X _13986_/B _13984_/Y _14350_/A vssd1 vssd1 vccd1 vccd1 _13985_/X
+ sky130_fd_sc_hd__o211a_1
X_16773_ _18042_/CLK _16773_/D vssd1 vssd1 vccd1 vccd1 _16773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15724_ _17730_/CLK _15724_/D vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _12936_/A _12936_/B vssd1 vssd1 vccd1 vccd1 _17488_/D sky130_fd_sc_hd__and2_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18443_ _18454_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _17262_/CLK _15655_/D vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfxtp_1
X_12867_ _12924_/A _12867_/B vssd1 vssd1 vccd1 vccd1 _17465_/D sky130_fd_sc_hd__and2_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _15215_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__nand2_1
X_11818_ hold4871/X _13811_/B _11817_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _11818_/X
+ sky130_fd_sc_hd__o211a_1
X_18374_ _18420_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
X_15586_ _17718_/CLK _15586_/D vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12798_ _12825_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _17442_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_248_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17274_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17528_/CLK hold347/X vssd1 vssd1 vccd1 vccd1 _17325_/Q sky130_fd_sc_hd__dfxtp_1
X_14537_ _15217_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14537_/Y sky130_fd_sc_hd__nand2_1
X_11749_ _12331_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_172_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17256_ _17453_/CLK _17256_/D vssd1 vssd1 vccd1 vccd1 _17256_/Q sky130_fd_sc_hd__dfxtp_1
X_14468_ hold2538/X _14481_/B _14467_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ _13710_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13419_/X sky130_fd_sc_hd__or2_1
X_16207_ _17439_/CLK _16207_/D vssd1 vssd1 vccd1 vccd1 _16207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17187_ _17283_/CLK _17187_/D vssd1 vssd1 vccd1 vccd1 _17187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _14740_/A _14411_/B vssd1 vssd1 vccd1 vccd1 _14399_/X sky130_fd_sc_hd__or2_1
X_16138_ _17313_/CLK _16138_/D vssd1 vssd1 vccd1 vccd1 hold512/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08960_ _15454_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _16097_/D sky130_fd_sc_hd__and2_1
X_16069_ _17287_/CLK _16069_/D vssd1 vssd1 vccd1 vccd1 hold650/A sky130_fd_sc_hd__dfxtp_1
Xhold3207 _10171_/X vssd1 vssd1 vccd1 vccd1 _16547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3218 _13321_/X vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3229 _12917_/X vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__dlygate4sd3_1
X_07911_ hold2106/X _07918_/B _07910_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _07911_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2506 _14013_/X vssd1 vssd1 vccd1 vccd1 _17812_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08891_ _15344_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__and2_1
Xhold2517 _07951_/X vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2528 _15677_/Q vssd1 vssd1 vccd1 vccd1 hold2528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 _14468_/X vssd1 vssd1 vccd1 vccd1 _18031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _14564_/X vssd1 vssd1 vccd1 vccd1 hold1805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 _15630_/Q vssd1 vssd1 vccd1 vccd1 hold1816/X sky130_fd_sc_hd__dlygate4sd3_1
X_07842_ hold2399/X _07865_/B _07841_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _07842_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1827 _07981_/X vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1838 _15885_/Q vssd1 vssd1 vccd1 vccd1 hold1838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1849 _17992_/Q vssd1 vssd1 vccd1 vccd1 hold1849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ _18241_/Q _13094_/A _11153_/C vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ _09447_/C _09447_/D _09442_/Y vssd1 vssd1 vccd1 vccd1 _09443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ hold331/X _09365_/B _09362_/D hold591/X _09373_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ _15549_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _14529_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08187_ _14246_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08187_/X sky130_fd_sc_hd__or2_1
Xhold5110 _17651_/Q vssd1 vssd1 vccd1 vccd1 hold5110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5121 _09568_/X vssd1 vssd1 vccd1 vccd1 _16346_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5132 _17672_/Q vssd1 vssd1 vccd1 vccd1 hold5132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5143 _10462_/X vssd1 vssd1 vccd1 vccd1 _16644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5154 _16554_/Q vssd1 vssd1 vccd1 vccd1 hold5154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4420 _11452_/X vssd1 vssd1 vccd1 vccd1 _16974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5165 _13375_/X vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5176 _09781_/X vssd1 vssd1 vccd1 vccd1 _16417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4431 _16933_/Q vssd1 vssd1 vccd1 vccd1 hold4431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5187 _16417_/Q vssd1 vssd1 vccd1 vccd1 hold5187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4442 _11362_/X vssd1 vssd1 vccd1 vccd1 _16944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4453 _16575_/Q vssd1 vssd1 vccd1 vccd1 hold4453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5198 _10369_/X vssd1 vssd1 vccd1 vccd1 _16613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4464 _13543_/X vssd1 vssd1 vccd1 vccd1 _17634_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3730 _10642_/Y vssd1 vssd1 vccd1 vccd1 _16704_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4475 _16861_/Q vssd1 vssd1 vccd1 vccd1 hold4475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3741 _12376_/Y vssd1 vssd1 vccd1 vccd1 _17282_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10080_ _10380_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10080_/X sky130_fd_sc_hd__or2_1
Xhold4486 _17219_/Q vssd1 vssd1 vccd1 vccd1 hold4486/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4497 _13336_/X vssd1 vssd1 vccd1 vccd1 _17565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3752 _11145_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3763 _09631_/X vssd1 vssd1 vccd1 vccd1 _16367_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3774 _12316_/Y vssd1 vssd1 vccd1 vccd1 _17262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3785 _11187_/Y vssd1 vssd1 vccd1 vccd1 _11188_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3796 _17112_/Q vssd1 vssd1 vccd1 vccd1 hold3796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13770_ _13770_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__or2_1
X_10982_ hold2036/X _16818_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12721_ hold1898/X hold3511/X _12805_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ hold389/X _09365_/B _09362_/D hold294/X _15438_/X vssd1 vssd1 vccd1 vccd1
+ _15442_/C sky130_fd_sc_hd__a221o_1
X_12652_ hold1760/X hold3099/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ hold829/X _17025_/Q _12152_/S vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__mux2_1
X_15371_ _16301_/Q _15477_/A2 _15487_/B1 hold679/X _15370_/X vssd1 vssd1 vccd1 vccd1
+ _15372_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12583_ hold2123/X hold2302/X _12679_/S vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17110_ _17898_/CLK _17110_/D vssd1 vssd1 vccd1 vccd1 _17110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14322_ _15217_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__nand2_1
X_18090_ _18226_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
X_11534_ hold1881/X hold4205/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17041_ _17889_/CLK _17041_/D vssd1 vssd1 vccd1 vccd1 _17041_/Q sky130_fd_sc_hd__dfxtp_1
X_14253_ hold2899/X _14272_/B _14252_/X _15072_/A vssd1 vssd1 vccd1 vccd1 _14253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11465_ hold841/X _16979_/Q _11753_/C vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ hold3784/X _13203_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__mux2_1
X_10416_ _10542_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14184_ hold747/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14184_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ hold2328/X _16956_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ _13183_/A1 _13133_/X _13134_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _11103_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__or2_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _17559_/Q _17093_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__mux2_1
X_17943_ _18071_/CLK hold786/X vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_1
X_10278_ _10563_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12017_ hold2681/X _17163_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__mux2_1
X_17874_ _17898_/CLK hold588/X vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
X_16825_ _18208_/CLK _16825_/D vssd1 vssd1 vccd1 vccd1 _16825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16756_ _18055_/CLK _16756_/D vssd1 vssd1 vccd1 vccd1 _16756_/Q sky130_fd_sc_hd__dfxtp_1
X_13968_ _15529_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13968_/X sky130_fd_sc_hd__or2_1
X_15707_ _17275_/CLK _15707_/D vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ hold2767/X hold3265/X _12919_/S vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__mux2_1
X_16687_ _18218_/CLK _16687_/D vssd1 vssd1 vccd1 vccd1 _16687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ _14352_/A _13899_/B vssd1 vssd1 vccd1 vccd1 _17757_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18426_ _18426_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15638_ _17268_/CLK _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18389_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15569_ _17779_/CLK _15569_/D vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _14850_/A hold1442/X hold196/X vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__mux2_1
X_17308_ _18405_/CLK _17308_/D vssd1 vssd1 vccd1 vccd1 hold393/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09090_ _15531_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__or2_1
X_18288_ _18390_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08041_ _14728_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08041_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ _17907_/CLK _17239_/D vssd1 vssd1 vccd1 vccd1 _17239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold902 hold902/A vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold913 hold913/A vssd1 vssd1 vccd1 vccd1 hold913/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold924 becStatus[1] vssd1 vssd1 vccd1 vccd1 input2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold935 hold935/A vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold946 hold946/A vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3004 _17477_/Q vssd1 vssd1 vccd1 vccd1 hold3004/X sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _16488_/Q _09992_/B _11066_/S vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__and3_1
Xhold979 hold979/A vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3015 _12635_/X vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3026 _12752_/X vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ hold32/X hold679/X _08993_/S vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__mux2_1
Xhold3037 _17382_/Q vssd1 vssd1 vccd1 vccd1 hold3037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3048 _17438_/Q vssd1 vssd1 vccd1 vccd1 hold3048/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2303 _12587_/X vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2314 _16274_/Q vssd1 vssd1 vccd1 vccd1 hold2314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3059 _17499_/Q vssd1 vssd1 vccd1 vccd1 hold3059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 _14416_/X vssd1 vssd1 vccd1 vccd1 _18006_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2336 _15681_/Q vssd1 vssd1 vccd1 vccd1 hold2336/X sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ hold407/X hold454/X _08932_/S vssd1 vssd1 vccd1 vccd1 hold455/A sky130_fd_sc_hd__mux2_1
Xhold2347 _15230_/X vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _09439_/X vssd1 vssd1 vccd1 vccd1 _16305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 _14853_/X vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _15542_/X vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _09421_/X vssd1 vssd1 vccd1 vccd1 _16296_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _15825_/Q vssd1 vssd1 vccd1 vccd1 hold2369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 _08182_/X vssd1 vssd1 vccd1 vccd1 _15727_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 _16257_/Q vssd1 vssd1 vccd1 vccd1 hold1646/X sky130_fd_sc_hd__dlygate4sd3_1
X_07825_ _07809_/X _07810_/Y hold1773/X _15477_/A2 vssd1 vssd1 vccd1 vccd1 _07825_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _16288_/Q vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 _09075_/X vssd1 vssd1 vccd1 vccd1 _16152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 _17784_/Q vssd1 vssd1 vccd1 vccd1 hold1679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09426_ _09438_/B _16299_/Q vssd1 vssd1 vccd1 vccd1 _09426_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _09357_/A _09392_/A vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__or2_2
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08308_ hold1189/X _08323_/B _08307_/X _13723_/C1 vssd1 vssd1 vccd1 vccd1 _08308_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09288_ hold1067/X _09338_/A2 _09287_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08239_ hold1335/X _08268_/B _08238_/X _08345_/A vssd1 vssd1 vccd1 vccd1 _08239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _11637_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_127_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10201_ hold3334/X _10589_/B _10200_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10201_/X
+ sky130_fd_sc_hd__o211a_1
X_11181_ hold3849/X _11097_/A _11180_/X vssd1 vssd1 vccd1 vccd1 _11181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4250 _16819_/Q vssd1 vssd1 vccd1 vccd1 hold4250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4261 _17222_/Q vssd1 vssd1 vccd1 vccd1 hold4261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10132_ hold4542/X _10646_/B _10131_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _10132_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4272 _10300_/X vssd1 vssd1 vccd1 vccd1 _16590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4283 hold4720/X vssd1 vssd1 vccd1 vccd1 hold4283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4294 _09601_/X vssd1 vssd1 vccd1 vccd1 _16357_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3560 _17673_/Q vssd1 vssd1 vccd1 vccd1 hold3560/X sky130_fd_sc_hd__dlygate4sd3_1
X_10063_ _10588_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10063_/Y sky130_fd_sc_hd__nor2_1
Xhold3571 _13657_/X vssd1 vssd1 vccd1 vccd1 _17672_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14940_ _15209_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14940_/X sky130_fd_sc_hd__or2_1
Xhold3582 _12542_/X vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3593 _17490_/Q vssd1 vssd1 vccd1 vccd1 hold3593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2870 _15589_/Q vssd1 vssd1 vccd1 vccd1 hold2870/X sky130_fd_sc_hd__dlygate4sd3_1
X_14871_ hold1559/X _14880_/B _14870_/X _14889_/C1 vssd1 vssd1 vccd1 vccd1 _14871_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2881 _14651_/X vssd1 vssd1 vccd1 vccd1 _18118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2892 _14869_/X vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16610_ _18218_/CLK _16610_/D vssd1 vssd1 vccd1 vccd1 _16610_/Q sky130_fd_sc_hd__dfxtp_1
X_13822_ _13822_/A _13822_/B vssd1 vssd1 vccd1 vccd1 _13822_/Y sky130_fd_sc_hd__nor2_1
X_17590_ _17686_/CLK _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _18131_/CLK _16541_/D vssd1 vssd1 vccd1 vccd1 _16541_/Q sky130_fd_sc_hd__dfxtp_1
X_13753_ hold3482/X _13847_/B _13752_/X _13753_/C1 vssd1 vssd1 vccd1 vccd1 _13753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ _11061_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ hold3466/X _12703_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13684_ hold3564/X _13886_/B _13683_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _13684_/X
+ sky130_fd_sc_hd__o211a_1
X_16472_ _18353_/CLK _16472_/D vssd1 vssd1 vccd1 vccd1 _16472_/Q sky130_fd_sc_hd__dfxtp_1
X_10896_ _10998_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18211_ _18266_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
X_15423_ _15481_/A1 _15415_/X _15422_/X _15481_/B1 hold5865/A vssd1 vssd1 vccd1 vccd1
+ _15423_/X sky130_fd_sc_hd__a32o_1
X_12635_ hold3014/X _12634_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_128_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18142_ _18235_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
X_15354_ _15354_/A _15354_/B vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__and2_1
X_12566_ hold3590/X _12565_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__mux2_1
X_11517_ _12093_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__or2_1
X_14305_ hold2715/X _14333_/A2 _14304_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ hold506/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15285_/X sky130_fd_sc_hd__or2_1
X_18073_ _18073_/CLK hold852/X vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
X_12497_ hold50/X _12509_/A2 _12505_/A3 _12496_/X _09003_/A vssd1 vssd1 vccd1 vccd1
+ hold51/A sky130_fd_sc_hd__o311a_1
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17024_ _17904_/CLK _17024_/D vssd1 vssd1 vccd1 vccd1 _17024_/Q sky130_fd_sc_hd__dfxtp_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__buf_6
X_14236_ _14970_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _11640_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14167_ hold1138/X _14198_/B _14166_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _14167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _11667_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__or2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__or2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _15551_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14098_/X sky130_fd_sc_hd__or2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13046_/A _13053_/A _13055_/C vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _18208_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
X_17857_ _17923_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _18431_/CLK _16808_/D vssd1 vssd1 vccd1 vccd1 _16808_/Q sky130_fd_sc_hd__dfxtp_1
X_08590_ hold380/X hold645/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_263_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17788_ _18427_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16739_ _18069_/CLK _16739_/D vssd1 vssd1 vccd1 vccd1 _16739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09211_ hold1355/X _09218_/B _09210_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _09211_/X
+ sky130_fd_sc_hd__o211a_1
X_18409_ _18409_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09142_ _15525_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09073_ hold2628/X _09119_/A2 _09072_/X _12936_/A vssd1 vssd1 vccd1 vccd1 _09073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08024_ hold2295/X _08029_/B _08023_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _08024_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 hold721/A vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold732 hold732/A vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 hold888/X vssd1 vssd1 vccd1 vccd1 hold889/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold765 hold765/A vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 hold776/A vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 la_data_in[14] vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__or2_1
Xhold798 hold879/X vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2100 _18341_/Q vssd1 vssd1 vccd1 vccd1 hold2100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2111 _15738_/Q vssd1 vssd1 vccd1 vccd1 hold2111/X sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ hold359/X hold482/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__mux2_1
Xhold2122 _09177_/X vssd1 vssd1 vccd1 vccd1 _16201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _15638_/Q vssd1 vssd1 vccd1 vccd1 hold2133/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2144 _08099_/X vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _18354_/Q vssd1 vssd1 vccd1 vccd1 hold1410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 _18041_/Q vssd1 vssd1 vccd1 vccd1 hold2155/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2166 _09324_/X vssd1 vssd1 vccd1 vccd1 _16272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 _13014_/X vssd1 vssd1 vccd1 vccd1 _17515_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ _15050_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _16047_/D sky130_fd_sc_hd__and2_1
Xhold1432 _18250_/Q vssd1 vssd1 vccd1 vccd1 hold1432/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2177 hold2177/A vssd1 vssd1 vccd1 vccd1 _12836_/S sky130_fd_sc_hd__buf_6
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2188 _14649_/X vssd1 vssd1 vccd1 vccd1 _18117_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1443 _17956_/Q vssd1 vssd1 vccd1 vccd1 hold1443/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1454 _08312_/X vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2199 _15798_/Q vssd1 vssd1 vccd1 vccd1 hold2199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 _16164_/Q vssd1 vssd1 vccd1 vccd1 hold1465/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ _12442_/A _13048_/A hold1915/X _07807_/X vssd1 vssd1 vccd1 vccd1 _07808_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1476 _14277_/X vssd1 vssd1 vccd1 vccd1 _17939_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _15454_/A hold360/X vssd1 vssd1 vccd1 vccd1 _16014_/D sky130_fd_sc_hd__and2_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _15094_/X vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _08059_/X vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ hold4145/X _11735_/B _10749_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _10750_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ _07804_/A _09447_/B _15334_/A _09408_/X vssd1 vssd1 vccd1 vccd1 _09409_/X
+ sky130_fd_sc_hd__o211a_1
X_10681_ hold4605/X _11735_/B _10680_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _10681_/X
+ sky130_fd_sc_hd__o211a_1
X_12420_ _12420_/A _12420_/B vssd1 vssd1 vccd1 vccd1 _17303_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ hold3153/X _12279_/A _12350_/X vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_67_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17329_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11302_ hold5005/X _11741_/B _11301_/X _13933_/A vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__o211a_1
X_15070_ _15070_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__and2_1
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12282_ _12282_/A _12282_/B vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14021_ hold2607/X _14040_/B _14020_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14021_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ hold4431/X _11617_/A2 _11232_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11164_ _11203_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11164_/Y sky130_fd_sc_hd__nor2_1
Xhold4080 _10390_/X vssd1 vssd1 vccd1 vccd1 _16620_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10115_ hold2872/X _16529_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__mux2_1
Xhold4091 _16841_/Q vssd1 vssd1 vccd1 vccd1 hold4091/X sky130_fd_sc_hd__dlygate4sd3_1
X_15972_ _18407_/CLK _15972_/D vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__dfxtp_1
X_11095_ _11189_/A _11216_/B _11094_/X _14390_/A vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__o211a_1
X_17711_ _17743_/CLK _17711_/D vssd1 vssd1 vccd1 vccd1 _17711_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3390 _17611_/Q vssd1 vssd1 vccd1 vccd1 hold3390/X sky130_fd_sc_hd__dlygate4sd3_1
X_14923_ hold5948/X _14946_/B hold366/X _15364_/A vssd1 vssd1 vccd1 vccd1 hold367/A
+ sky130_fd_sc_hd__o211a_1
X_10046_ _16506_/Q _10070_/B _10271_/S vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__and3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__buf_4
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__buf_1
X_17642_ _17708_/CLK _17642_/D vssd1 vssd1 vccd1 vccd1 _17642_/Q sky130_fd_sc_hd__dfxtp_1
X_14854_ _14854_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__or2_1
X_13805_ _17722_/Q _13805_/B _13805_/C vssd1 vssd1 vccd1 vccd1 _13805_/X sky130_fd_sc_hd__and3_1
X_17573_ _17739_/CLK _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
X_14785_ hold2799/X _14772_/B _14784_/X _14881_/C1 vssd1 vssd1 vccd1 vccd1 _14785_/X
+ sky130_fd_sc_hd__o211a_1
X_11997_ _12093_/A _11997_/B vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16524_ _18210_/CLK _16524_/D vssd1 vssd1 vccd1 vccd1 _16524_/Q sky130_fd_sc_hd__dfxtp_1
X_13736_ hold985/X hold4345/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__mux2_1
X_10948_ hold3479/X _11732_/B _10947_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _10948_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16455_ _18304_/CLK _16455_/D vssd1 vssd1 vccd1 vccd1 _16455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13667_ hold1418/X _17676_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__mux2_1
X_10879_ hold5719/X _11201_/B _10878_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _17344_/Q _15486_/B1 _15485_/B1 hold372/X vssd1 vssd1 vccd1 vccd1 _15406_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _12885_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _17382_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16386_ _18395_/CLK _16386_/D vssd1 vssd1 vccd1 vccd1 _16386_/Q sky130_fd_sc_hd__dfxtp_1
X_13598_ _15786_/Q _17653_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13599_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18125_ _18197_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15337_ hold247/X _09357_/A _15484_/B1 hold447/X _15336_/X vssd1 vssd1 vccd1 vccd1
+ _15342_/B sky130_fd_sc_hd__a221o_1
X_12549_ _12924_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _17359_/D sky130_fd_sc_hd__and2_1
XFILLER_0_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5709 _16991_/Q vssd1 vssd1 vccd1 vccd1 hold5709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_1 _13197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056_ _18066_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
X_15268_ hold721/X _09386_/A _09392_/D hold594/X vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _17855_/CLK _17007_/D vssd1 vssd1 vccd1 vccd1 _17007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ hold1956/X _14216_/Y _14218_/X _14492_/C1 vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15199_ _15199_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 _10610_/C vssd1 vssd1 vccd1 vccd1 _10643_/C sky130_fd_sc_hd__clkbuf_8
Xfanout519 fanout523/X vssd1 vssd1 vccd1 vccd1 _10649_/C sky130_fd_sc_hd__buf_4
X_09760_ hold3548/X _10070_/B _09759_/X _15144_/C1 vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__o211a_1
X_08711_ hold149/X hold306/X _08727_/S vssd1 vssd1 vccd1 vccd1 _08712_/B sky130_fd_sc_hd__mux2_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _18427_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_1
X_09691_ hold5150/X _10073_/B _09690_/X _15030_/A vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08642_ _15304_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _15943_/D sky130_fd_sc_hd__and2_1
XFILLER_0_117_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08573_ _12430_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _15910_/D sky130_fd_sc_hd__and2_1
XFILLER_0_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ hold607/X _15508_/B vssd1 vssd1 vccd1 vccd1 _09170_/B sky130_fd_sc_hd__or2_2
X_09056_ hold359/X hold713/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08007_ _15521_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08007_/X sky130_fd_sc_hd__or2_1
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__buf_4
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold551 hold551/A vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 hold562/A vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold573/A vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__buf_6
Xhold584 data_in[30] vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 hold595/A vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ hold4573/X _10070_/B _09957_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09958_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_185_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18118_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _12422_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _16072_/D sky130_fd_sc_hd__and2_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ hold5664/X _10016_/B _09888_/X _15060_/A vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18337_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1240 _15875_/Q vssd1 vssd1 vccd1 vccd1 hold1240/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 _15624_/Q vssd1 vssd1 vccd1 vccd1 hold1251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1262 _08475_/X vssd1 vssd1 vccd1 vccd1 _15866_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ hold4218/X _13811_/B _11919_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _11920_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1273 _15594_/Q vssd1 vssd1 vccd1 vccd1 hold1273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 _15587_/Q vssd1 vssd1 vccd1 vccd1 hold1284/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _14410_/X vssd1 vssd1 vccd1 vccd1 _18003_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ hold5348/X _12329_/B _11850_/X _13931_/A vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ hold2304/X hold4591/X _11192_/C vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__mux2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _15492_/A _14573_/B hold1813/X vssd1 vssd1 vccd1 vccd1 _14570_/X sky130_fd_sc_hd__a21o_1
X_11782_ _12331_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _11782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _13710_/A _13521_/B vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__or2_1
X_10733_ hold2080/X hold5266/X _11213_/C vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13452_ _13776_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__or2_1
X_16240_ _17428_/CLK _16240_/D vssd1 vssd1 vccd1 vccd1 _16240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ hold1461/X hold3751/X _11732_/C vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12403_ hold136/X hold561/X _12443_/S vssd1 vssd1 vccd1 vccd1 hold562/A sky130_fd_sc_hd__mux2_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13383_ _13674_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_1
X_16171_ _17517_/CLK _16171_/D vssd1 vssd1 vccd1 vccd1 _16171_/Q sky130_fd_sc_hd__dfxtp_1
X_10595_ _10595_/A _10619_/B _10619_/C vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ _13873_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__nor2_1
X_15122_ hold2135/X _15109_/B _15121_/X _15168_/C1 vssd1 vssd1 vccd1 vccd1 _15122_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ hold265/X _18312_/Q hold302/A vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ hold4953/X _13871_/B _12264_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _12265_/X
+ sky130_fd_sc_hd__o211a_1
X_14004_ hold756/X _14052_/B vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ _16896_/Q _11216_/B _11216_/C vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__and3_1
X_12196_ hold4267/X _12308_/B _12195_/X _08161_/A vssd1 vssd1 vccd1 vccd1 _12196_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput82 _13209_/A vssd1 vssd1 vccd1 vccd1 output82/X sky130_fd_sc_hd__buf_6
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 _13289_/A vssd1 vssd1 vccd1 vccd1 output93/X sky130_fd_sc_hd__buf_6
X_11147_ _16873_/Q _11150_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__and3_1
XFILLER_0_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15955_ _17302_/CLK _15955_/D vssd1 vssd1 vccd1 vccd1 hold550/A sky130_fd_sc_hd__dfxtp_1
X_11078_ hold2992/X hold4228/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10029_ _13190_/A _09933_/A _10028_/X vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__a21oi_1
X_14906_ hold490/X _14910_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or2_1
X_15886_ _17724_/CLK _15886_/D vssd1 vssd1 vccd1 vccd1 _15886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17625_ _17721_/CLK _17625_/D vssd1 vssd1 vccd1 vccd1 _17625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ hold2603/X _14828_/B _14836_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14837_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _18223_/CLK _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14768_ _15000_/A _14774_/B vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16507_ _18396_/CLK _16507_/D vssd1 vssd1 vccd1 vccd1 _16507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _13800_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13719_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17487_ _17487_/CLK _17487_/D vssd1 vssd1 vccd1 vccd1 _17487_/Q sky130_fd_sc_hd__dfxtp_1
X_14699_ hold2930/X _14720_/B _14698_/X _14831_/C1 vssd1 vssd1 vccd1 vccd1 _14699_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16438_ _18383_/CLK _16438_/D vssd1 vssd1 vccd1 vccd1 _16438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16369_ _18378_/CLK _16369_/D vssd1 vssd1 vccd1 vccd1 _16369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18108_ _18205_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5506 _17086_/Q vssd1 vssd1 vccd1 vccd1 hold5506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5517 _09613_/X vssd1 vssd1 vccd1 vccd1 _16361_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5528 _16454_/Q vssd1 vssd1 vccd1 vccd1 hold5528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5539 _11023_/X vssd1 vssd1 vccd1 vccd1 _16831_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4805 _17627_/Q vssd1 vssd1 vccd1 vccd1 hold4805/X sky130_fd_sc_hd__dlygate4sd3_1
X_18039_ _18305_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
Xhold4816 _17648_/Q vssd1 vssd1 vccd1 vccd1 hold4816/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4827 _13459_/X vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4838 _17669_/Q vssd1 vssd1 vccd1 vccd1 hold4838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4849 _13678_/X vssd1 vssd1 vccd1 vccd1 _17679_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _09981_/A vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout316 _10560_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__buf_4
Xfanout327 fanout337/X vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__buf_2
X_09812_ hold2100/X _16428_/Q _10010_/C vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__mux2_1
Xfanout338 _12508_/B vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__buf_4
Xfanout349 _08965_/S vssd1 vssd1 vccd1 vccd1 _08997_/S sky130_fd_sc_hd__buf_8
X_09743_ hold2117/X hold3283/X _10010_/C vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09674_ hold2433/X _16382_/Q _10562_/S vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08625_ hold59/X hold611/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08626_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ hold81/X hold557/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__mux2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08487_ hold875/X _08486_/B _08486_/Y _08133_/A vssd1 vssd1 vccd1 vccd1 hold876/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ _15169_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__or2_1
X_09039_ _15284_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _16136_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ hold2441/X hold5397/X _12338_/C vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__mux2_1
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold381 hold381/A vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 hold392/A vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _11103_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout850 _11203_/A vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__buf_6
XFILLER_0_102_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout861 _07785_/Y vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__buf_4
XFILLER_0_99_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout872 _15221_/A vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__clkbuf_16
Xfanout883 hold967/X vssd1 vssd1 vccd1 vccd1 hold949/A sky130_fd_sc_hd__buf_6
Xfanout894 hold490/X vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__buf_8
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _17743_/CLK _15740_/D vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ hold2858/X hold3572/X _12955_/S vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__mux2_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 hold1070/A vssd1 vssd1 vccd1 vccd1 input53/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _16239_/Q vssd1 vssd1 vccd1 vccd1 hold1081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ hold2397/X hold4379/X _13796_/S vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__mux2_1
Xhold1092 _15106_/X vssd1 vssd1 vccd1 vccd1 _18337_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _18428_/CLK _15671_/D vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ hold2599/X _17472_/Q _12910_/S vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux2_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17439_/CLK _17410_/D vssd1 vssd1 vccd1 vccd1 _17410_/Q sky130_fd_sc_hd__dfxtp_1
X_14622_ _15231_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14622_/X sky130_fd_sc_hd__or2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18390_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
X_11834_ hold1442/X _17102_/Q _12353_/C vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/CLK hold51/X vssd1 vssd1 vccd1 vccd1 _17341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11765_ _17079_/Q _11765_/B _11765_/C vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__and3_1
X_14553_ hold784/X _14553_/B vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_leaf_84_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17340_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ hold3526/X _13880_/B _13503_/X _13792_/C1 vssd1 vssd1 vccd1 vccd1 _13504_/X
+ sky130_fd_sc_hd__o211a_1
X_10716_ _11667_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__or2_1
X_17272_ _17282_/CLK _17272_/D vssd1 vssd1 vccd1 vccd1 _17272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18454_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11696_ hold2270/X _17056_/Q _11792_/C vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__mux2_1
X_14484_ hold1790/X _14487_/B _14483_/Y _15044_/A vssd1 vssd1 vccd1 vccd1 _14484_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16223_ _17456_/CLK _16223_/D vssd1 vssd1 vccd1 vccd1 _16223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ hold3699/X _10521_/A _10646_/X vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__a21oi_1
X_13435_ hold3422/X _13862_/B _13434_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ hold5086/X _13844_/B _13365_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _13366_/X
+ sky130_fd_sc_hd__o211a_1
X_16154_ _17494_/CLK _16154_/D vssd1 vssd1 vccd1 vccd1 _16154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ hold3144/X _10098_/A _10577_/X vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15105_ _15105_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15105_/X sky130_fd_sc_hd__or2_1
X_12317_ _17263_/Q _12356_/B _12356_/C vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__and3_1
X_13297_ _13297_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13297_/X sky130_fd_sc_hd__and2_1
X_16085_ _17284_/CLK _16085_/D vssd1 vssd1 vccd1 vccd1 hold456/A sky130_fd_sc_hd__dfxtp_1
X_12248_ hold1370/X hold4862/X _13844_/C vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__mux2_1
X_15036_ _15036_/A hold950/X vssd1 vssd1 vccd1 vccd1 hold951/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ hold2168/X _17217_/Q _13844_/C vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16987_ _17855_/CLK _16987_/D vssd1 vssd1 vccd1 vccd1 _16987_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _17289_/CLK _15938_/D vssd1 vssd1 vccd1 vccd1 hold409/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15869_ _17736_/CLK _15869_/D vssd1 vssd1 vccd1 vccd1 _15869_/Q sky130_fd_sc_hd__dfxtp_1
X_08410_ hold1187/X _08440_/A2 _08409_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _08410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17608_ _17738_/CLK _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_1
X_09390_ _09369_/C _09389_/X _18460_/Q vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _08389_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _15802_/D sky130_fd_sc_hd__and2_1
X_17539_ _18386_/CLK _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ _15551_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08272_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6004 _18416_/Q vssd1 vssd1 vccd1 vccd1 hold6004/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6015 data_in[3] vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6026 _16326_/Q vssd1 vssd1 vccd1 vccd1 hold6026/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6037 _17525_/Q vssd1 vssd1 vccd1 vccd1 hold6037/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5303 _16338_/Q vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5314 _11164_/Y vssd1 vssd1 vccd1 vccd1 _16878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5325 _11763_/Y vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5336 _16494_/Q vssd1 vssd1 vccd1 vccd1 hold5336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4602 _11590_/X vssd1 vssd1 vccd1 vccd1 _17020_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5347 _10903_/X vssd1 vssd1 vccd1 vccd1 _16791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5358 _11770_/Y vssd1 vssd1 vccd1 vccd1 _17080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4613 _17069_/Q vssd1 vssd1 vccd1 vccd1 hold4613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4624 _12013_/X vssd1 vssd1 vccd1 vccd1 _17161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5369 _17203_/Q vssd1 vssd1 vccd1 vccd1 hold5369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4635 _17283_/Q vssd1 vssd1 vccd1 vccd1 hold4635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3901 _10047_/Y vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4646 _11086_/X vssd1 vssd1 vccd1 vccd1 _16852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4657 _16560_/Q vssd1 vssd1 vccd1 vccd1 hold4657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3912 _16519_/Q vssd1 vssd1 vccd1 vccd1 hold3912/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4668 _12274_/X vssd1 vssd1 vccd1 vccd1 _17248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3923 _10822_/X vssd1 vssd1 vccd1 vccd1 _16764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3934 _15997_/Q vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4679 _16686_/Q vssd1 vssd1 vccd1 vccd1 hold4679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3945 _17584_/Q vssd1 vssd1 vccd1 vccd1 hold3945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3956 _15333_/X vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3967 _16702_/Q vssd1 vssd1 vccd1 vccd1 hold3967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3978 _16892_/Q vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold3989 hold5831/X vssd1 vssd1 vccd1 vccd1 hold3989/X sky130_fd_sc_hd__clkbuf_4
Xfanout157 _12836_/S vssd1 vssd1 vccd1 vccd1 _12980_/S sky130_fd_sc_hd__buf_6
Xfanout168 _09494_/X vssd1 vssd1 vccd1 vccd1 _13823_/B sky130_fd_sc_hd__buf_2
X_07987_ hold2689/X _07991_/A2 _07986_/X _13411_/C1 vssd1 vssd1 vccd1 vccd1 _07987_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout179 _10852_/A2 vssd1 vssd1 vccd1 vccd1 _11741_/B sky130_fd_sc_hd__clkbuf_4
X_09726_ _09918_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__or2_1
X_09657_ _11082_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _12430_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _15926_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09951_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__or2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _12420_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _15893_/D sky130_fd_sc_hd__and2_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ _12036_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11550_/X sky130_fd_sc_hd__or2_1
X_10501_ _10595_/A _10619_/B _10500_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _16657_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _12153_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ hold3708/X _13219_/X _13300_/S vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__mux2_1
X_10432_ hold3305/X _10640_/B _10431_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ _13183_/A1 _13149_/X _13150_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13151_/X
+ sky130_fd_sc_hd__o211a_1
X_10363_ hold4151/X _10640_/B _10362_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _12210_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5870 _18423_/Q vssd1 vssd1 vccd1 vccd1 hold5870/X sky130_fd_sc_hd__dlygate4sd3_1
X_13082_ _17561_/Q _17095_/Q _13250_/S vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__mux2_1
Xhold5881 _18463_/X vssd1 vssd1 vccd1 vccd1 hold5881/X sky130_fd_sc_hd__buf_1
X_10294_ hold4155/X _10580_/B _10293_/X _14807_/C1 vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5892 _07794_/Y vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12033_ _13794_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__or2_1
X_16910_ _18051_/CLK _16910_/D vssd1 vssd1 vccd1 vccd1 _16910_/Q sky130_fd_sc_hd__dfxtp_1
X_17890_ _17890_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _18013_/CLK _16841_/D vssd1 vssd1 vccd1 vccd1 _16841_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout680 _14418_/C1 vssd1 vssd1 vccd1 vccd1 _14492_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout691 _15244_/A vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__buf_2
X_16772_ _18071_/CLK _16772_/D vssd1 vssd1 vccd1 vccd1 _16772_/Q sky130_fd_sc_hd__dfxtp_1
X_13984_ _15545_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15723_ _17257_/CLK _15723_/D vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ hold3042/X _12934_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__mux2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _18451_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _17262_/CLK _15654_/D vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12866_ hold3289/X _12865_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__mux2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ hold1161/X _14612_/B _14604_/X _14887_/C1 vssd1 vssd1 vccd1 vccd1 _14605_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18373_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
X_11817_ _13716_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__or2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15585_ _17253_/CLK _15585_/D vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ hold3119/X _12796_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17524_/CLK hold127/X vssd1 vssd1 vccd1 vccd1 _17324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ hold2386/X _14541_/B _14535_/Y _13935_/A vssd1 vssd1 vccd1 vccd1 _14536_/X
+ sky130_fd_sc_hd__o211a_1
X_11748_ hold3645/X _11652_/A _11747_/X vssd1 vssd1 vccd1 vccd1 _11748_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17255_ _17453_/CLK _17255_/D vssd1 vssd1 vccd1 vccd1 _17255_/Q sky130_fd_sc_hd__dfxtp_1
X_14467_ _14986_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14467_/X sky130_fd_sc_hd__or2_1
X_11679_ _11688_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_288_wb_clk_i clkbuf_5_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16206_ _17439_/CLK _16206_/D vssd1 vssd1 vccd1 vccd1 _16206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ hold2961/X _17593_/Q _13805_/C vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17186_ _17703_/CLK _17186_/D vssd1 vssd1 vccd1 vccd1 _17186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ hold1300/X hold209/X _14397_/X _14392_/A vssd1 vssd1 vccd1 vccd1 _14398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_217_wb_clk_i clkbuf_5_23__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16137_ _17331_/CLK _16137_/D vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ hold2435/X _17570_/Q _13829_/C vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16068_ _18406_/CLK _16068_/D vssd1 vssd1 vccd1 vccd1 hold568/A sky130_fd_sc_hd__dfxtp_1
Xhold3208 _16836_/Q vssd1 vssd1 vccd1 vccd1 hold3208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3219 _16599_/Q vssd1 vssd1 vccd1 vccd1 hold3219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07910_ _15533_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__or2_1
X_15019_ hold2433/X _15006_/B _15018_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _15019_/X
+ sky130_fd_sc_hd__o211a_1
X_08890_ hold53/X hold311/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__mux2_1
Xhold2507 _18216_/Q vssd1 vssd1 vccd1 vccd1 hold2507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 _18399_/Q vssd1 vssd1 vccd1 vccd1 hold2518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 _08075_/X vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07841_ _14854_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__or2_1
Xhold1806 _14565_/X vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1817 _07975_/X vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 _15886_/Q vssd1 vssd1 vccd1 vccd1 hold1828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 _08516_/X vssd1 vssd1 vccd1 vccd1 _15885_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09511_ hold5592/X _09998_/B _09510_/X _15394_/A vssd1 vssd1 vccd1 vccd1 _09511_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ _09447_/C _09447_/D _09481_/B vssd1 vssd1 vccd1 vccd1 _09442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _17325_/Q _09357_/A _09392_/B hold722/X vssd1 vssd1 vccd1 vccd1 _09373_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ hold1820/X _08336_/A2 _08323_/Y _09272_/A vssd1 vssd1 vccd1 vccd1 _08324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08255_ hold2588/X _08262_/B _08254_/X _08349_/A vssd1 vssd1 vccd1 vccd1 _08255_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ hold2411/X _08209_/B _08185_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _08186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5100 _16381_/Q vssd1 vssd1 vccd1 vccd1 hold5100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5111 _13498_/X vssd1 vssd1 vccd1 vccd1 _17619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5122 _17609_/Q vssd1 vssd1 vccd1 vccd1 hold5122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5133 _13561_/X vssd1 vssd1 vccd1 vccd1 _17640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5144 _17705_/Q vssd1 vssd1 vccd1 vccd1 hold5144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4410 _11698_/X vssd1 vssd1 vccd1 vccd1 _17056_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5155 _10096_/X vssd1 vssd1 vccd1 vccd1 _16522_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5166 _16008_/Q vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4421 _16324_/Q vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__buf_1
Xhold5177 _17706_/Q vssd1 vssd1 vccd1 vccd1 hold5177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4432 _11233_/X vssd1 vssd1 vccd1 vccd1 _16901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4443 _17223_/Q vssd1 vssd1 vccd1 vccd1 hold4443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5188 _09685_/X vssd1 vssd1 vccd1 vccd1 _16385_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4454 _10159_/X vssd1 vssd1 vccd1 vccd1 _16543_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5199 hold5838/X vssd1 vssd1 vccd1 vccd1 hold5839/A sky130_fd_sc_hd__buf_4
Xhold4465 _17633_/Q vssd1 vssd1 vccd1 vccd1 hold4465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3720 _11727_/Y vssd1 vssd1 vccd1 vccd1 _11728_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3731 _17118_/Q vssd1 vssd1 vccd1 vccd1 hold3731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4476 _11017_/X vssd1 vssd1 vccd1 vccd1 _16829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4487 _12091_/X vssd1 vssd1 vccd1 vccd1 _17187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3742 _16909_/Q vssd1 vssd1 vccd1 vccd1 hold3742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4498 _17614_/Q vssd1 vssd1 vccd1 vccd1 hold4498/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3753 _11146_/Y vssd1 vssd1 vccd1 vccd1 _16872_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3764 _17566_/Q vssd1 vssd1 vccd1 vccd1 hold3764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3775 _17096_/Q vssd1 vssd1 vccd1 vccd1 hold3775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3786 _11188_/Y vssd1 vssd1 vccd1 vccd1 _16886_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3797 _12345_/Y vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__dlygate4sd3_1
X_09709_ hold5641/X _09998_/B _09708_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__o211a_1
X_10981_ hold3299/X _11171_/B _10980_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _10981_/X
+ sky130_fd_sc_hd__o211a_1
X_12720_ _12813_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _17416_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ _12825_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _17393_/D sky130_fd_sc_hd__and2_1
XFILLER_0_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ hold4694/X _11792_/B _11601_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__o211a_1
X_15370_ hold435/X _15486_/A2 _15446_/B1 hold563/X vssd1 vssd1 vccd1 vccd1 _15370_/X
+ sky130_fd_sc_hd__a22o_1
X_12582_ _12987_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _17370_/D sky130_fd_sc_hd__and2_1
XFILLER_0_33_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ hold1002/X _14326_/B _14320_/Y _14733_/C1 vssd1 vssd1 vccd1 vccd1 _14321_/X
+ sky130_fd_sc_hd__o211a_1
X_11533_ hold4391/X _11726_/B _11532_/X _15504_/A vssd1 vssd1 vccd1 vccd1 _11533_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ _17856_/CLK _17040_/D vssd1 vssd1 vccd1 vccd1 _17040_/Q sky130_fd_sc_hd__dfxtp_1
X_11464_ hold5460/X _11753_/B _11463_/X _14380_/A vssd1 vssd1 vccd1 vccd1 _11464_/X
+ sky130_fd_sc_hd__o211a_1
X_14252_ _14986_/A _14280_/B vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_310_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _18187_/Q hold4051/X _10637_/C vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__mux2_1
X_13203_ _13202_/X _16918_/Q _13307_/S vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__mux2_1
X_11395_ hold4508/X _12320_/B _11394_/X _14193_/C1 vssd1 vssd1 vccd1 vccd1 _11395_/X
+ sky130_fd_sc_hd__o211a_1
X_14183_ hold1084/X _14202_/B _14182_/X _14191_/C1 vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__o211a_1
X_13134_ _13134_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__or2_1
X_10346_ hold2897/X _16606_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__mux2_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__and2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _18003_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
X_10277_ hold2930/X _16583_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__mux2_1
X_12016_ hold4343/X _13811_/B _12015_/X _08355_/A vssd1 vssd1 vccd1 vccd1 _12016_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17873_ _17873_/CLK hold830/X vssd1 vssd1 vccd1 vccd1 hold829/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16824_ _18059_/CLK _16824_/D vssd1 vssd1 vccd1 vccd1 _16824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16755_ _18208_/CLK _16755_/D vssd1 vssd1 vccd1 vccd1 _16755_/Q sky130_fd_sc_hd__dfxtp_1
X_13967_ hold2417/X _13980_/B _13966_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__o211a_1
X_15706_ _17703_/CLK _15706_/D vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _12918_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _17482_/D sky130_fd_sc_hd__and2_1
X_16686_ _18265_/CLK _16686_/D vssd1 vssd1 vccd1 vccd1 _16686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _15513_/A hold2886/X hold244/X vssd1 vssd1 vccd1 vccd1 _13899_/B sky130_fd_sc_hd__mux2_1
X_18425_ _18425_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15637_ _17266_/CLK _15637_/D vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12849_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _17459_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18356_ _18390_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15568_ _17268_/CLK _15568_/D vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17307_ _17307_/CLK _17307_/D vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
X_14519_ _14984_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__or2_1
XFILLER_0_142_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18287_ _18319_/CLK hold868/X vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15499_ _15515_/A hold1584/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15500_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ hold1983/X _08033_/B _08039_/X _08147_/A vssd1 vssd1 vccd1 vccd1 _08040_/X
+ sky130_fd_sc_hd__o211a_1
X_17238_ _17906_/CLK _17238_/D vssd1 vssd1 vccd1 vccd1 _17238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold914 hold914/A vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _17902_/CLK _17169_/D vssd1 vssd1 vccd1 vccd1 _17169_/Q sky130_fd_sc_hd__dfxtp_1
Xhold925 input2/X vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold936 hold936/A vssd1 vssd1 vccd1 vccd1 hold936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold947 hold964/X vssd1 vssd1 vccd1 vccd1 hold965/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _11155_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3005 _12902_/X vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3016 _17402_/Q vssd1 vssd1 vccd1 vccd1 hold3016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3027 _17426_/Q vssd1 vssd1 vccd1 vccd1 hold3027/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08942_ _09063_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _16088_/D sky130_fd_sc_hd__and2_1
Xhold3038 _17423_/Q vssd1 vssd1 vccd1 vccd1 hold3038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3049 _12785_/X vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2304 _17961_/Q vssd1 vssd1 vccd1 vccd1 hold2304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _09328_/X vssd1 vssd1 vccd1 vccd1 _16274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _15687_/Q vssd1 vssd1 vccd1 vccd1 hold2326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2337 _08083_/X vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08873_ _12430_/A hold386/X vssd1 vssd1 vccd1 vccd1 _16054_/D sky130_fd_sc_hd__and2_1
Xhold1603 _15704_/Q vssd1 vssd1 vccd1 vccd1 hold1603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _16198_/Q vssd1 vssd1 vccd1 vccd1 hold2348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1614 _18297_/Q vssd1 vssd1 vccd1 vccd1 hold1614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 _18126_/Q vssd1 vssd1 vccd1 vccd1 hold2359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1625 _17810_/Q vssd1 vssd1 vccd1 vccd1 hold1625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1636 hold6038/X vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__buf_1
X_07824_ _09400_/A _09122_/A _07824_/C _09121_/B vssd1 vssd1 vccd1 vccd1 _07824_/Y
+ sky130_fd_sc_hd__nor4_2
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1647 _09294_/X vssd1 vssd1 vccd1 vccd1 _16257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 _09405_/X vssd1 vssd1 vccd1 vccd1 _16288_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 _15805_/Q vssd1 vssd1 vccd1 vccd1 hold1669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ _07804_/A _09472_/C _15304_/A _09424_/X vssd1 vssd1 vccd1 vccd1 _09425_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09356_ _09400_/A _09366_/B _09356_/C vssd1 vssd1 vccd1 vccd1 _09356_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_75_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_139_wb_clk_i clkbuf_5_27__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18388_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _15531_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08307_/X sky130_fd_sc_hd__or2_1
X_09287_ _15183_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ _14511_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _08171_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__and2_1
X_10200_ _10527_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__or2_1
XFILLER_0_160_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ _16884_/Q _11192_/B _11192_/C vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4240 _16573_/Q vssd1 vssd1 vccd1 vccd1 hold4240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4251 _10891_/X vssd1 vssd1 vccd1 vccd1 _16787_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10131_ _10521_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__or2_1
Xhold4262 _12100_/X vssd1 vssd1 vccd1 vccd1 _17190_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4273 _16574_/Q vssd1 vssd1 vccd1 vccd1 hold4273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4284 _13735_/X vssd1 vssd1 vccd1 vccd1 _17698_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3550 _17641_/Q vssd1 vssd1 vccd1 vccd1 hold3550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4295 _16568_/Q vssd1 vssd1 vccd1 vccd1 hold4295/X sky130_fd_sc_hd__dlygate4sd3_1
X_10062_ _13278_/A _10506_/A _10061_/X vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__a21oi_1
Xhold3561 _13564_/X vssd1 vssd1 vccd1 vccd1 _17641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3572 _17495_/Q vssd1 vssd1 vccd1 vccd1 hold3572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3583 _17494_/Q vssd1 vssd1 vccd1 vccd1 hold3583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3594 _17358_/Q vssd1 vssd1 vccd1 vccd1 hold3594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2860 _15641_/Q vssd1 vssd1 vccd1 vccd1 hold2860/X sky130_fd_sc_hd__dlygate4sd3_1
X_14870_ _15209_/A _14894_/B vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__or2_1
Xhold2871 _07891_/X vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2882 _18107_/Q vssd1 vssd1 vccd1 vccd1 hold2882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 _18084_/Q vssd1 vssd1 vccd1 vccd1 hold2893/X sky130_fd_sc_hd__dlygate4sd3_1
X_13821_ hold3687/X _13734_/A _13820_/X vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _18206_/CLK _16540_/D vssd1 vssd1 vccd1 vccd1 _16540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _13758_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10964_ hold2094/X hold3985/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ hold997/X hold3384/X _12820_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _18392_/CLK _16471_/D vssd1 vssd1 vccd1 vccd1 _16471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13683_ _13779_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ hold1849/X _16789_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_183_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _18210_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
X_15422_ _15471_/A _15422_/B _15422_/C _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/X
+ sky130_fd_sc_hd__or4_1
X_12634_ hold1014/X _17389_/Q _12676_/S vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _18205_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15353_ _15481_/A1 _15345_/X _15352_/X _15481_/B1 hold5185/X vssd1 vssd1 vccd1 vccd1
+ _15353_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12565_ hold2370/X _17366_/Q _12955_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ _14984_/A _14338_/B vssd1 vssd1 vccd1 vccd1 _14304_/X sky130_fd_sc_hd__or2_1
XFILLER_0_145_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ hold1265/X hold3442/X _12320_/C vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__mux2_1
X_18072_ _18072_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
X_15284_ _15284_/A _15284_/B vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__and2_1
X_12496_ _17341_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17023_ _17903_/CLK _17023_/D vssd1 vssd1 vccd1 vccd1 _17023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14235_ hold1016/X _14266_/B _14234_/X _15044_/A vssd1 vssd1 vccd1 vccd1 _14235_/X
+ sky130_fd_sc_hd__o211a_1
X_11447_ hold2147/X _16973_/Q _11735_/C vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14166_ hold892/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14166_/X sky130_fd_sc_hd__or2_1
X_11378_ hold975/X _16950_/Q _11762_/C vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__mux2_1
X_13117_ _13116_/X hold3144/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10998_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__or2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ hold1896/X _14094_/B _14096_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14097_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13048_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__and2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _18053_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_1
X_17856_ _17856_/CLK hold880/X vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _17981_/CLK _16807_/D vssd1 vssd1 vccd1 vccd1 _16807_/Q sky130_fd_sc_hd__dfxtp_1
X_17787_ _17852_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
X_14999_ hold1385/X _15004_/B _14998_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _14999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ _18032_/CLK _16738_/D vssd1 vssd1 vccd1 vccd1 _16738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16669_ _18227_/CLK _16669_/D vssd1 vssd1 vccd1 vccd1 _16669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _15539_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__or2_1
X_18408_ _18408_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_232_wb_clk_i clkbuf_5_21__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17205_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09141_ hold1073/X _09177_/A2 _09140_/X _12876_/A vssd1 vssd1 vccd1 vccd1 _09141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18339_ _18339_/CLK hold864/X vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ _14972_/A _09118_/B vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08023_ _15537_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08023_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 hold700/A vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold711 hold711/A vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 hold722/A vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold733 hold787/X vssd1 vssd1 vccd1 vccd1 hold788/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 hold744/A vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 hold890/X vssd1 vssd1 vccd1 vccd1 hold891/A sky130_fd_sc_hd__buf_6
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 la_data_in[22] vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 hold788/A vssd1 vssd1 vccd1 vccd1 input42/A sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ hold1718/X hold4753/X _10271_/S vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__mux2_1
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__buf_8
Xhold2101 _15114_/X vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2112 _08204_/X vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08925_ _15284_/A _08925_/B vssd1 vssd1 vccd1 vccd1 _16080_/D sky130_fd_sc_hd__and2_1
Xhold2123 _16270_/Q vssd1 vssd1 vccd1 vccd1 hold2123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2134 _07991_/X vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2145 _15664_/Q vssd1 vssd1 vccd1 vccd1 hold2145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 _14452_/X vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1411 _15142_/X vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 _14488_/X vssd1 vssd1 vccd1 vccd1 _18041_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1422 _15582_/Q vssd1 vssd1 vccd1 vccd1 hold1422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 _17984_/Q vssd1 vssd1 vccd1 vccd1 hold2167/X sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ hold65/X hold117/X _08864_/S vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__mux2_1
Xhold1433 _14927_/X vssd1 vssd1 vccd1 vccd1 _18250_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2178 _12644_/X vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 _15679_/Q vssd1 vssd1 vccd1 vccd1 hold2189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 _14313_/X vssd1 vssd1 vccd1 vccd1 _17956_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1455 _15686_/Q vssd1 vssd1 vccd1 vccd1 hold1455/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1466 _09099_/X vssd1 vssd1 vccd1 vccd1 _16164_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ _07785_/Y _18462_/Q _07805_/A _07806_/Y vssd1 vssd1 vccd1 vccd1 _07807_/X
+ sky130_fd_sc_hd__a22o_1
Xhold1477 _18317_/Q vssd1 vssd1 vccd1 vccd1 hold1477/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08787_ hold359/X _16014_/Q _08787_/S vssd1 vssd1 vccd1 vccd1 hold360/A sky130_fd_sc_hd__mux2_1
Xhold1488 _17991_/Q vssd1 vssd1 vccd1 vccd1 hold1488/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _18212_/Q vssd1 vssd1 vccd1 vccd1 hold1499/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _09438_/B _16290_/Q vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__or2_1
X_10680_ _11640_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09339_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _17274_/Q _12374_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__and3_1
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _12036_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12281_ hold1885/X _17251_/Q _12377_/C vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11232_ _12018_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11232_/X sky130_fd_sc_hd__or2_1
X_14020_ _15527_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11163_ hold5312/X _11106_/A _11162_/X vssd1 vssd1 vccd1 vccd1 _11163_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_wb_clk_i clkbuf_5_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18071_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4070 _13507_/X vssd1 vssd1 vccd1 vccd1 _17622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4081 _16380_/Q vssd1 vssd1 vccd1 vccd1 hold4081/X sky130_fd_sc_hd__dlygate4sd3_1
X_10114_ hold4657/X _10568_/B _10113_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10114_/X
+ sky130_fd_sc_hd__o211a_1
X_15971_ _18410_/CLK _15971_/D vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11094_ _11121_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11094_/X sky130_fd_sc_hd__or2_1
Xhold4092 _10957_/X vssd1 vssd1 vccd1 vccd1 _16809_/D sky130_fd_sc_hd__dlygate4sd3_1
X_17710_ _17742_/CLK _17710_/D vssd1 vssd1 vccd1 vccd1 _17710_/Q sky130_fd_sc_hd__dfxtp_1
Xhold3380 _17492_/Q vssd1 vssd1 vccd1 vccd1 hold3380/X sky130_fd_sc_hd__dlygate4sd3_1
X_10045_ _10588_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10045_/Y sky130_fd_sc_hd__nor2_1
X_14922_ hold490/A _14964_/B vssd1 vssd1 vccd1 vccd1 hold366/A sky130_fd_sc_hd__or2_1
Xhold3391 _13378_/X vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__clkbuf_4
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _17649_/CLK _17641_/D vssd1 vssd1 vccd1 vccd1 _17641_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2690 _07987_/X vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ hold1612/X _14880_/B _14852_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14853_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ _13822_/A _13804_/B vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17572_ _17739_/CLK _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
X_14784_ _15231_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14784_/X sky130_fd_sc_hd__or2_1
X_11996_ hold2522/X _17156_/Q _12320_/C vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16523_ _18392_/CLK _16523_/D vssd1 vssd1 vccd1 vccd1 _16523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ _13829_/A _13829_/B _13734_/X _08367_/A vssd1 vssd1 vccd1 vccd1 _13735_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10947_ _11616_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16454_ _18337_/CLK _16454_/D vssd1 vssd1 vccd1 vccd1 _16454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ hold4969/X _13856_/B _13665_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13666_/X
+ sky130_fd_sc_hd__o211a_1
X_10878_ _11106_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10878_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15405_ _15405_/A _15483_/B vssd1 vssd1 vccd1 vccd1 _15405_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ hold3037/X _12616_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__mux2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _18330_/CLK _16385_/D vssd1 vssd1 vccd1 vccd1 _16385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ hold5207/X _13883_/B _13596_/X _08391_/A vssd1 vssd1 vccd1 vccd1 _13597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18124_ _18140_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
X_15336_ _17337_/Q _09362_/C _15485_/B1 hold453/X vssd1 vssd1 vccd1 vccd1 _15336_/X
+ sky130_fd_sc_hd__a22o_1
X_12548_ hold3236/X _12547_/X _12926_/S vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ _18055_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ hold724/X _15479_/A2 _09386_/D hold520/X _15266_/X vssd1 vssd1 vccd1 vccd1
+ _15272_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12479_ hold20/X _08598_/B _08999_/B _12478_/X _09047_/A vssd1 vssd1 vccd1 vccd1
+ hold21/A sky130_fd_sc_hd__o311a_1
XANTENNA_2 _13197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17006_ _18051_/CLK _17006_/D vssd1 vssd1 vccd1 vccd1 _17006_/Q sky130_fd_sc_hd__dfxtp_1
X_14218_ _14218_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14218_/X sky130_fd_sc_hd__or2_1
X_15198_ hold1540/X _15219_/B _15197_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14149_ hold2060/X _14148_/B _14148_/Y _14149_/C1 vssd1 vssd1 vccd1 vccd1 _14149_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout509 _10610_/C vssd1 vssd1 vccd1 vccd1 _10625_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08710_ _15394_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__and2_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _17908_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_1
X_09690_ _10506_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__or2_1
X_08641_ hold8/X hold592/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__mux2_1
X_17839_ _17903_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_5_19__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_19__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_08572_ hold5/X hold138/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ hold607/X _15508_/B vssd1 vssd1 vccd1 vccd1 _09124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ _12420_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _16144_/D sky130_fd_sc_hd__and2_1
XFILLER_0_170_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ hold2522/X _08029_/B _08005_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _08006_/X
+ sky130_fd_sc_hd__o211a_1
Xhold530 hold530/A vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 hold552/A vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold563 hold563/A vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 hold574/A vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__buf_2
Xhold596 hold596/A vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ _09975_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__or2_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ hold17/X hold371/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__mux2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09987_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__or2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _13951_/X vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _08493_/X vssd1 vssd1 vccd1 vccd1 _15875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 _07963_/X vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ _15344_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _16038_/D sky130_fd_sc_hd__and2_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1263 _16180_/Q vssd1 vssd1 vccd1 vccd1 hold1263/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1274 _07901_/X vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _07887_/X vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 la_data_in[2] vssd1 vssd1 vccd1 vccd1 hold1296/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _12234_/A _11850_/B vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__or2_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_154_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ hold5391/X _10897_/A2 _10800_/X _14344_/A vssd1 vssd1 vccd1 vccd1 _10801_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ hold3799/X _12036_/A _11780_/X vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ hold1843/X _17627_/Q _13805_/C vssd1 vssd1 vccd1 vccd1 _13521_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10732_ hold5594/X _11762_/B _10731_/X _13917_/A vssd1 vssd1 vccd1 vccd1 _10732_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13451_ hold1716/X hold4480/X _13868_/C vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ hold5413/X _11150_/B _10662_/X _14368_/A vssd1 vssd1 vccd1 vccd1 _10663_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _12402_/A _12402_/B vssd1 vssd1 vccd1 vccd1 _17294_/D sky130_fd_sc_hd__and2_1
X_16170_ _17506_/CLK _16170_/D vssd1 vssd1 vccd1 vccd1 _16170_/Q sky130_fd_sc_hd__dfxtp_1
X_10594_ _11194_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10594_/Y sky130_fd_sc_hd__nor2_1
X_13382_ hold2006/X hold3138/X _13832_/C vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__mux2_1
X_15121_ _15229_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__or2_1
X_12333_ hold3174/X _12243_/A _12332_/X vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15052_ _15052_/A hold981/X vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__and2_1
X_12264_ _13392_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14003_ hold1357/X _14036_/B _14002_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _14003_/X
+ sky130_fd_sc_hd__o211a_1
X_11215_ _11218_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _11215_/Y sky130_fd_sc_hd__nor2_1
X_12195_ _13797_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput72 _13051_/A vssd1 vssd1 vccd1 vccd1 output72/X sky130_fd_sc_hd__buf_6
Xoutput83 _13065_/A vssd1 vssd1 vccd1 vccd1 output83/X sky130_fd_sc_hd__buf_6
X_11146_ _12301_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 _13073_/A vssd1 vssd1 vccd1 vccd1 output94/X sky130_fd_sc_hd__buf_6
X_15954_ _17307_/CLK _15954_/D vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__dfxtp_1
X_11077_ hold3373/X _11171_/B _11076_/X _13901_/A vssd1 vssd1 vccd1 vccd1 _11077_/X
+ sky130_fd_sc_hd__o211a_1
X_10028_ _16500_/Q _10028_/B _10028_/C vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__and3_1
X_14905_ hold5954/X hold657/A hold638/X _14905_/C1 vssd1 vssd1 vccd1 vccd1 hold639/A
+ sky130_fd_sc_hd__o211a_1
X_15885_ _17722_/CLK _15885_/D vssd1 vssd1 vccd1 vccd1 _15885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17624_ _17725_/CLK _17624_/D vssd1 vssd1 vccd1 vccd1 _17624_/Q sky130_fd_sc_hd__dfxtp_1
X_14836_ _15229_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14836_/X sky130_fd_sc_hd__or2_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17555_ _18229_/CLK _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14767_ hold1469/X _14772_/B _14766_/X _14875_/C1 vssd1 vssd1 vccd1 vccd1 _14767_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _13392_/A _11979_/B vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16506_ _18396_/CLK _16506_/D vssd1 vssd1 vccd1 vccd1 _16506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13718_ hold2568/X hold4226/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__mux2_1
X_17486_ _17494_/CLK _17486_/D vssd1 vssd1 vccd1 vccd1 _17486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14698_ _14984_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ _18381_/CLK _16437_/D vssd1 vssd1 vccd1 vccd1 _16437_/Q sky130_fd_sc_hd__dfxtp_1
X_13649_ hold1022/X _17670_/Q _13859_/C vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16368_ _18391_/CLK _16368_/D vssd1 vssd1 vccd1 vccd1 _16368_/Q sky130_fd_sc_hd__dfxtp_1
X_18107_ _18267_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_1
X_15319_ hold221/X _15485_/A2 _15447_/B1 hold307/X _15318_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5507 _11692_/X vssd1 vssd1 vccd1 vccd1 _17054_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16299_ _18460_/CLK _16299_/D vssd1 vssd1 vccd1 vccd1 _16299_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5518 _16800_/Q vssd1 vssd1 vccd1 vccd1 hold5518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5529 _09796_/X vssd1 vssd1 vccd1 vccd1 _16422_/D sky130_fd_sc_hd__dlygate4sd3_1
X_18038_ _18070_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4806 _13426_/X vssd1 vssd1 vccd1 vccd1 _17595_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4817 _13489_/X vssd1 vssd1 vccd1 vccd1 _17616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4828 _17596_/Q vssd1 vssd1 vccd1 vccd1 hold4828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4839 _13552_/X vssd1 vssd1 vccd1 vccd1 _17637_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout306 _09981_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_4
X_09811_ hold3833/X _10001_/B _09810_/X _14985_/C1 vssd1 vssd1 vccd1 vccd1 _09811_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout317 fanout337/X vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__buf_2
Xfanout328 _10098_/A vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__buf_4
Xfanout339 _12506_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__buf_4
X_09742_ hold3263/X _10013_/B _09741_/X _15064_/A vssd1 vssd1 vccd1 vccd1 _09742_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ hold4467/X _10049_/B _09672_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09673_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08970_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _15934_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _12422_/A hold340/X vssd1 vssd1 vccd1 vccd1 _15901_/D sky130_fd_sc_hd__and2_1
X_08486_ _14950_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ hold762/X _09106_/B _09106_/Y _12984_/A vssd1 vssd1 vccd1 vccd1 hold763/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ hold17/X hold98/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold360 hold360/A vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold382/A vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 hold393/A vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ hold2985/X hold5550/X _11213_/C vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__mux2_1
Xfanout840 fanout841/X vssd1 vssd1 vccd1 vccd1 _14865_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout851 _11791_/A vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__buf_8
Xfanout862 _15215_/A vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__buf_12
Xfanout873 _07780_/Y vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__buf_12
Xfanout884 _15195_/A vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__buf_8
XFILLER_0_99_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 hold667/X vssd1 vssd1 vccd1 vccd1 _15515_/A sky130_fd_sc_hd__buf_8
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _17493_/D sky130_fd_sc_hd__and2_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1060 _14795_/X vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 input53/X vssd1 vssd1 vccd1 vccd1 hold1071/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ hold5162/X _12305_/B _11901_/X _15498_/A vssd1 vssd1 vccd1 vccd1 _11902_/X
+ sky130_fd_sc_hd__o211a_1
X_15670_ _17221_/CLK _15670_/D vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1082 _17840_/Q vssd1 vssd1 vccd1 vccd1 hold1082/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _15813_/Q vssd1 vssd1 vccd1 vccd1 hold1093/X sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _12885_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _17470_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ hold2592/X _14612_/B _14620_/X _14867_/C1 vssd1 vssd1 vccd1 vccd1 _14621_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ hold5042/X _12311_/B _11832_/X _08109_/A vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17340_ _17340_/CLK hold189/X vssd1 vssd1 vccd1 vccd1 _17340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ hold2969/X _14554_/A2 _14551_/X _13897_/A vssd1 vssd1 vccd1 vccd1 _14552_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _12343_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13503_ _13791_/A _13503_/B vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__or2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17907_/CLK _17271_/D vssd1 vssd1 vccd1 vccd1 _17271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ hold2308/X hold5263/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_126_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14483_ _15543_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__nand2_1
X_11695_ hold5713/X _11789_/B _11694_/X _13935_/A vssd1 vssd1 vccd1 vccd1 _11695_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16222_ _17453_/CLK _16222_/D vssd1 vssd1 vccd1 vccd1 _16222_/Q sky130_fd_sc_hd__dfxtp_1
X_13434_ _13734_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _13434_/X sky130_fd_sc_hd__or2_1
X_10646_ _16706_/Q _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16153_ _17506_/CLK _16153_/D vssd1 vssd1 vccd1 vccd1 _16153_/Q sky130_fd_sc_hd__dfxtp_1
X_13365_ _13749_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__or2_1
X_10577_ _16683_/Q _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10577_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_51_wb_clk_i clkbuf_5_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ hold2159/X _15113_/B _15103_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _15104_/X
+ sky130_fd_sc_hd__o211a_1
X_12316_ _13822_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12316_/Y sky130_fd_sc_hd__nor2_1
X_16084_ _17329_/CLK _16084_/D vssd1 vssd1 vccd1 vccd1 hold394/A sky130_fd_sc_hd__dfxtp_1
X_13296_ _13289_/X _13295_/X _13304_/B1 vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15035_ hold949/X _18303_/Q hold302/X vssd1 vssd1 vccd1 vccd1 hold950/A sky130_fd_sc_hd__mux2_1
X_12247_ hold4923/X _12341_/B _12246_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__o211a_1
X_12178_ hold4733/X _12377_/B _12177_/X _12274_/C1 vssd1 vssd1 vccd1 vccd1 _12178_/X
+ sky130_fd_sc_hd__o211a_1
X_11129_ hold1911/X _16867_/Q _11765_/C vssd1 vssd1 vccd1 vccd1 _11130_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _17896_/CLK _16986_/D vssd1 vssd1 vccd1 vccd1 _16986_/Q sky130_fd_sc_hd__dfxtp_1
X_15937_ _17284_/CLK _15937_/D vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _17739_/CLK hold809/X vssd1 vssd1 vccd1 vccd1 hold808/A sky130_fd_sc_hd__dfxtp_1
X_17607_ _17735_/CLK _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_1
X_14819_ hold2226/X _14828_/B _14818_/X _14885_/C1 vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15799_ _17666_/CLK _15799_/D vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08340_ hold944/X hold1503/X hold122/X vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__mux2_1
X_17538_ _18386_/CLK _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ hold1987/X _08268_/B _08270_/X _08359_/A vssd1 vssd1 vccd1 vccd1 _08271_/X
+ sky130_fd_sc_hd__o211a_1
X_17469_ _17482_/CLK _17469_/D vssd1 vssd1 vccd1 vccd1 _17469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6005 _18420_/Q vssd1 vssd1 vccd1 vccd1 hold6005/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold6016 data_in[5] vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6027 la_data_in[3] vssd1 vssd1 vccd1 vccd1 hold664/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6038 _16311_/Q vssd1 vssd1 vccd1 vccd1 hold6038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5304 _10023_/Y vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5315 _16336_/Q vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5326 _11764_/Y vssd1 vssd1 vccd1 vccd1 _17078_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5337 _09916_/X vssd1 vssd1 vccd1 vccd1 _16462_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5348 _17139_/Q vssd1 vssd1 vccd1 vccd1 hold5348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4603 _16940_/Q vssd1 vssd1 vccd1 vccd1 hold4603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5359 _16441_/Q vssd1 vssd1 vccd1 vccd1 hold5359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4614 _11641_/X vssd1 vssd1 vccd1 vccd1 _17037_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4625 _16765_/Q vssd1 vssd1 vccd1 vccd1 hold4625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4636 _12283_/X vssd1 vssd1 vccd1 vccd1 _17251_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3902 _17575_/Q vssd1 vssd1 vccd1 vccd1 hold3902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4647 _17026_/Q vssd1 vssd1 vccd1 vccd1 hold4647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3913 _10566_/Y vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4658 _10114_/X vssd1 vssd1 vccd1 vccd1 _16528_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4669 _17269_/Q vssd1 vssd1 vccd1 vccd1 hold4669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3924 _16664_/Q vssd1 vssd1 vccd1 vccd1 hold3924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3935 _15283_/X vssd1 vssd1 vccd1 vccd1 _15284_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3946 _13872_/Y vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3957 _16505_/Q vssd1 vssd1 vccd1 vccd1 hold3957/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout147 _12800_/S vssd1 vssd1 vccd1 vccd1 _12821_/S sky130_fd_sc_hd__buf_6
Xhold3968 _10540_/X vssd1 vssd1 vccd1 vccd1 _16670_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3979 _11110_/X vssd1 vssd1 vccd1 vccd1 _16860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout158 hold2176/X vssd1 vssd1 vccd1 vccd1 hold2177/A sky130_fd_sc_hd__buf_6
X_07986_ hold800/X _07988_/B vssd1 vssd1 vccd1 vccd1 _07986_/X sky130_fd_sc_hd__or2_1
Xfanout169 _12314_/B vssd1 vssd1 vccd1 vccd1 _12311_/B sky130_fd_sc_hd__buf_4
XFILLER_0_129_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09725_ _18312_/Q hold3762/X _10028_/C vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__mux2_1
X_09656_ hold835/X _16376_/Q _11177_/C vssd1 vssd1 vccd1 vccd1 _09657_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08607_ hold32/X hold419/X _08655_/S vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_145_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09587_ hold2118/X _13294_/A _10067_/C vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__mux2_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ hold35/X hold505/X _08594_/S vssd1 vssd1 vccd1 vccd1 _08539_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08469_ hold1280/X _08486_/B _08468_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08469_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ _10524_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ hold2163/X hold4514/X _12152_/S vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_162_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10431_ _10527_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _13150_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__or2_1
X_10362_ _10554_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__or2_1
X_12101_ hold2310/X hold3340/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__mux2_1
Xhold5860 hold5943/X vssd1 vssd1 vccd1 vccd1 hold5860/X sky130_fd_sc_hd__buf_2
XFILLER_0_104_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _13081_/A fanout2/X vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__and2_1
X_10293_ _10548_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__or2_1
Xhold5871 hold5871/A vssd1 vssd1 vccd1 vccd1 hold5871/X sky130_fd_sc_hd__clkbuf_4
Xhold5882 hold5936/X vssd1 vssd1 vccd1 vccd1 _17754_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5893 _16908_/Q vssd1 vssd1 vccd1 vccd1 hold5893/X sky130_fd_sc_hd__dlygate4sd3_1
X_12032_ hold2064/X hold4803/X _13793_/S vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__mux2_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _17884_/CLK _16840_/D vssd1 vssd1 vccd1 vccd1 _16840_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout670 _08137_/A vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__buf_4
Xfanout681 _14171_/C1 vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__buf_4
X_16771_ _18069_/CLK _16771_/D vssd1 vssd1 vccd1 vccd1 _16771_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout692 _15244_/A vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__clkbuf_4
X_13983_ hold975/X _13986_/B _13982_/Y _13917_/A vssd1 vssd1 vccd1 vccd1 hold976/A
+ sky130_fd_sc_hd__o211a_1
X_15722_ _17878_/CLK _15722_/D vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ hold1667/X _17489_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__mux2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15653_ _17252_/CLK _15653_/D vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfxtp_1
X_18441_ _18441_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ hold2586/X _17466_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__mux2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _15105_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14604_/X sky130_fd_sc_hd__or2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18380_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
X_11816_ hold1174/X hold3775/X _13811_/C vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15584_ _17252_/CLK _15584_/D vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ hold2662/X hold3087/X _12814_/S vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17323_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _17323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _15000_/A _14541_/B vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _17073_/Q _11747_/B _11747_/C vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__and3_1
XFILLER_0_172_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17254_ _17719_/CLK _17254_/D vssd1 vssd1 vccd1 vccd1 _17254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ hold2738/X _14487_/B _14465_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _14466_/X
+ sky130_fd_sc_hd__o211a_1
X_11678_ hold1750/X hold4113/X _11783_/C vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16205_ _17439_/CLK _16205_/D vssd1 vssd1 vccd1 vccd1 _16205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13417_ hold4135/X _13808_/B _13416_/X _13801_/C1 vssd1 vssd1 vccd1 vccd1 _13417_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10629_ hold4003/X _10563_/A _10628_/X vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__a21oi_1
X_17185_ _17217_/CLK _17185_/D vssd1 vssd1 vccd1 vccd1 _17185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14397_ hold756/X _14445_/B vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16136_ _17331_/CLK _16136_/D vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ hold4281/X _13832_/B _13347_/X _08371_/A vssd1 vssd1 vccd1 vccd1 _13348_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16067_ _17287_/CLK _16067_/D vssd1 vssd1 vccd1 vccd1 hold647/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _13311_/A1 _13277_/X _13278_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13279_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3209 _10942_/X vssd1 vssd1 vccd1 vccd1 _16804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_257_wb_clk_i clkbuf_5_16__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17669_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15018_ _15233_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__or2_1
Xhold2508 _14855_/X vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 _15234_/X vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ hold1008/X _07865_/B _07839_/X _08111_/A vssd1 vssd1 vccd1 vccd1 _07840_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1807 _15769_/Q vssd1 vssd1 vccd1 vccd1 hold1807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1818 _17876_/Q vssd1 vssd1 vccd1 vccd1 hold1818/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1829 _08518_/X vssd1 vssd1 vccd1 vccd1 _15886_/D sky130_fd_sc_hd__dlygate4sd3_1
X_16969_ _17882_/CLK _16969_/D vssd1 vssd1 vccd1 vccd1 _16969_/Q sky130_fd_sc_hd__dfxtp_1
X_09510_ _09903_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__or2_1
X_09441_ _09447_/D _09481_/B vssd1 vssd1 vccd1 vccd1 _16306_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _07805_/A _09362_/A _09386_/A hold672/X vssd1 vssd1 vccd1 vccd1 _09375_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _15547_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08254_ _15533_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08254_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08185_ _14854_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__or2_1
Xhold5101 _09577_/X vssd1 vssd1 vccd1 vccd1 _16349_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5112 _17181_/Q vssd1 vssd1 vccd1 vccd1 hold5112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5123 _13372_/X vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5134 _16387_/Q vssd1 vssd1 vccd1 vccd1 hold5134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5145 _13660_/X vssd1 vssd1 vccd1 vccd1 _17673_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4400 _11605_/X vssd1 vssd1 vccd1 vccd1 _17025_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4411 _17726_/Q vssd1 vssd1 vccd1 vccd1 hold4411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5156 _17708_/Q vssd1 vssd1 vccd1 vccd1 hold5156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5167 _15393_/X vssd1 vssd1 vccd1 vccd1 _15394_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4422 _09982_/X vssd1 vssd1 vccd1 vccd1 _16484_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5178 _13663_/X vssd1 vssd1 vccd1 vccd1 _17674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4433 _17258_/Q vssd1 vssd1 vccd1 vccd1 hold4433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5189 _16480_/Q vssd1 vssd1 vccd1 vccd1 hold5189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4444 _12103_/X vssd1 vssd1 vccd1 vccd1 _17191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4455 _16937_/Q vssd1 vssd1 vccd1 vccd1 hold4455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3710 _11194_/Y vssd1 vssd1 vccd1 vccd1 _16888_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4466 _13444_/X vssd1 vssd1 vccd1 vccd1 _17601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3721 _11728_/Y vssd1 vssd1 vccd1 vccd1 _17066_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3732 _12363_/Y vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4477 _17089_/Q vssd1 vssd1 vccd1 vccd1 hold4477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3743 _11736_/Y vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4488 _16813_/Q vssd1 vssd1 vccd1 vccd1 hold4488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3754 _16537_/Q vssd1 vssd1 vccd1 vccd1 hold3754/X sky130_fd_sc_hd__buf_1
Xhold4499 _13387_/X vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3765 _13818_/Y vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3776 _12297_/Y vssd1 vssd1 vccd1 vccd1 _12298_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3787 _16905_/Q vssd1 vssd1 vccd1 vccd1 hold3787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3798 _12346_/Y vssd1 vssd1 vccd1 vccd1 _17272_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07969_ hold2310/X _07978_/B _07968_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _07969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _09903_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__or2_1
X_10980_ _11076_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09639_ _09987_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ hold3093/X _12649_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _11697_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_167_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ hold3071/X _12580_/X _12980_/S vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _15215_/A _14326_/B vssd1 vssd1 vccd1 vccd1 _14320_/Y sky130_fd_sc_hd__nand2_1
X_11532_ _11631_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__or2_1
XFILLER_0_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ hold2940/X _14266_/B _14250_/X _15007_/C1 vssd1 vssd1 vccd1 vccd1 _14251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _11658_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _17576_/Q _17110_/Q _13306_/S vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__mux2_1
X_10414_ hold4299/X _10649_/B _10413_/X _14859_/C1 vssd1 vssd1 vccd1 vccd1 _10414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14182_ hold883/X _14214_/B vssd1 vssd1 vccd1 vccd1 _14182_/X sky130_fd_sc_hd__or2_1
X_11394_ _11649_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13133_ _13132_/X hold3852/X _13173_/S vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ hold4327/X _10631_/B _10344_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10345_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5690 _11668_/X vssd1 vssd1 vccd1 vccd1 _17046_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13064_ _13051_/X _13063_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17526_/D sky130_fd_sc_hd__o21a_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _18032_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_1
X_10276_ hold4735/X _10568_/B _10275_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _10276_/X
+ sky130_fd_sc_hd__o211a_1
X_12015_ _13716_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_178_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17872_ _17904_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16823_ _18067_/CLK _16823_/D vssd1 vssd1 vccd1 vccd1 _16823_/Q sky130_fd_sc_hd__dfxtp_1
X_13966_ _14986_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13966_/X sky130_fd_sc_hd__or2_1
X_16754_ _18053_/CLK _16754_/D vssd1 vssd1 vccd1 vccd1 _16754_/Q sky130_fd_sc_hd__dfxtp_1
X_15705_ _17583_/CLK _15705_/D vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfxtp_1
X_12917_ hold3228/X _12916_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__mux2_1
X_16685_ _18266_/CLK _16685_/D vssd1 vssd1 vccd1 vccd1 _16685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13897_ _13897_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _17756_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18424_ _18424_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12848_ hold3067/X _12847_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__mux2_1
X_15636_ _17232_/CLK _15636_/D vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18355_ _18355_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
X_15567_ _17865_/CLK _15567_/D vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfxtp_1
X_12779_ hold3448/X _12778_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12779_/X sky130_fd_sc_hd__mux2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ _17342_/CLK _17306_/D vssd1 vssd1 vccd1 vccd1 hold710/A sky130_fd_sc_hd__dfxtp_1
X_14518_ hold1424/X _14541_/B _14517_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14518_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18286_ _18382_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__and2_1
XFILLER_0_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17237_ _17779_/CLK _17237_/D vssd1 vssd1 vccd1 vccd1 _17237_/Q sky130_fd_sc_hd__dfxtp_1
X_14449_ _15129_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17168_ _17232_/CLK _17168_/D vssd1 vssd1 vccd1 vccd1 _17168_/Q sky130_fd_sc_hd__dfxtp_1
Xhold904 hold904/A vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 hold915/A vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 hold926/A vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold937 hold937/A vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ _17342_/CLK _16119_/D vssd1 vssd1 vccd1 vccd1 hold674/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 hold966/X vssd1 vssd1 vccd1 vccd1 hold967/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ _13086_/A _09903_/A _09989_/X vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__a21oi_1
X_17099_ _18428_/CLK _17099_/D vssd1 vssd1 vccd1 vccd1 _17099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3006 _17480_/Q vssd1 vssd1 vccd1 vccd1 hold3006/X sky130_fd_sc_hd__dlygate4sd3_1
X_08941_ hold35/X hold515/X _08997_/S vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__mux2_1
Xhold3017 _12677_/X vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3028 _12749_/X vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3039 _12740_/X vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2305 _14323_/X vssd1 vssd1 vccd1 vccd1 _17961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 _15609_/Q vssd1 vssd1 vccd1 vccd1 hold2316/X sky130_fd_sc_hd__dlygate4sd3_1
X_08872_ hold68/X _16054_/Q _08930_/S vssd1 vssd1 vccd1 vccd1 hold386/A sky130_fd_sc_hd__mux2_1
Xhold2327 _08095_/X vssd1 vssd1 vccd1 vccd1 _15687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 _18010_/Q vssd1 vssd1 vccd1 vccd1 hold2338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _15745_/Q vssd1 vssd1 vccd1 vccd1 hold1604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 _09171_/X vssd1 vssd1 vccd1 vccd1 _16198_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1615 _18146_/Q vssd1 vssd1 vccd1 vccd1 hold1615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 _14009_/X vssd1 vssd1 vccd1 vccd1 _17810_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07823_ hold235/X hold265/X _09496_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _09121_/B
+ sky130_fd_sc_hd__or4b_1
Xhold1637 _09415_/X vssd1 vssd1 vccd1 vccd1 _16293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _16265_/Q vssd1 vssd1 vccd1 vccd1 hold1648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 _18256_/Q vssd1 vssd1 vccd1 vccd1 hold1659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ _09438_/B _16298_/Q vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _15547_/A _15219_/A _09359_/C vssd1 vssd1 vccd1 vccd1 _09356_/C sky130_fd_sc_hd__or3_1
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ hold5980/X _08336_/A2 _08305_/X _08349_/A vssd1 vssd1 vccd1 vccd1 hold817/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09286_ _14913_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__or2_2
XFILLER_0_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08237_ hold1738/X _08262_/B _08236_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_wb_clk_i clkbuf_5_28__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18034_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08168_ _15519_/A hold2550/X _08170_/S vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_wb_clk_i clkbuf_leaf_40_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18415_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08099_ hold2143/X _08088_/B _08098_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _08099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4230 _17664_/Q vssd1 vssd1 vccd1 vccd1 hold4230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4241 _10153_/X vssd1 vssd1 vccd1 vccd1 _16541_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10130_ hold2884/X hold3135/X _10646_/C vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__mux2_1
Xhold4252 _16687_/Q vssd1 vssd1 vccd1 vccd1 hold4252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4263 _16694_/Q vssd1 vssd1 vccd1 vccd1 hold4263/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4274 _10156_/X vssd1 vssd1 vccd1 vccd1 _16542_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4285 _16634_/Q vssd1 vssd1 vccd1 vccd1 hold4285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3540 _13696_/X vssd1 vssd1 vccd1 vccd1 _17685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10061_ _10061_/A _10601_/B _10481_/S vssd1 vssd1 vccd1 vccd1 _10061_/X sky130_fd_sc_hd__and3_1
Xhold3551 _13468_/X vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4296 _10138_/X vssd1 vssd1 vccd1 vccd1 _16536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3562 _16375_/Q vssd1 vssd1 vccd1 vccd1 hold3562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3573 _17681_/Q vssd1 vssd1 vccd1 vccd1 hold3573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3584 _17486_/Q vssd1 vssd1 vccd1 vccd1 hold3584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2850 _17761_/Q vssd1 vssd1 vccd1 vccd1 hold2850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3595 _17366_/Q vssd1 vssd1 vccd1 vccd1 hold3595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2861 _08000_/X vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2872 _18087_/Q vssd1 vssd1 vccd1 vccd1 hold2872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2883 _14629_/X vssd1 vssd1 vccd1 vccd1 _18107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2894 _14581_/X vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13820_ _17727_/Q _13829_/B _13829_/C vssd1 vssd1 vccd1 vccd1 _13820_/X sky130_fd_sc_hd__and3_1
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ hold2791/X _17704_/Q _13847_/C vssd1 vssd1 vccd1 vccd1 _13752_/B sky130_fd_sc_hd__mux2_1
X_10963_ hold5570/X _11156_/B _10962_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10963_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _12789_/A _12702_/B vssd1 vssd1 vccd1 vccd1 _17410_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16470_ _18385_/CLK _16470_/D vssd1 vssd1 vccd1 vccd1 _16470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13682_ hold2588/X _17681_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__mux2_1
X_10894_ hold4757/X _11192_/B _10893_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _10894_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15421_ _17302_/Q _15451_/A2 _09386_/D hold558/X _15416_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_155_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ _12855_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _17387_/D sky130_fd_sc_hd__and2_1
XFILLER_0_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15352_ _15471_/A _15352_/B _15352_/C _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__or4_1
X_18140_ _18140_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
X_12564_ _12933_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _17364_/D sky130_fd_sc_hd__and2_1
X_14303_ hold1542/X _14333_/A2 _14302_/X _14362_/A vssd1 vssd1 vccd1 vccd1 _14303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ hold5007/X _12341_/B _11514_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _11515_/X
+ sky130_fd_sc_hd__o211a_1
X_18071_ _18071_/CLK hold921/X vssd1 vssd1 vccd1 vccd1 hold920/A sky130_fd_sc_hd__dfxtp_1
X_15283_ _15490_/A1 _15275_/X _15282_/X _15490_/B1 _18404_/Q vssd1 vssd1 vccd1 vccd1
+ _15283_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ hold251/A _08598_/B _12445_/B _12494_/X _15454_/A vssd1 vssd1 vccd1 vccd1
+ hold189/A sky130_fd_sc_hd__o311a_1
XFILLER_0_151_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _17870_/CLK _17022_/D vssd1 vssd1 vccd1 vccd1 _17022_/Q sky130_fd_sc_hd__dfxtp_1
X_14234_ _15183_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14234_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ hold4879/X _11617_/A2 _11445_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _11446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ hold2732/X _14198_/B _14164_/X _14352_/A vssd1 vssd1 vccd1 vccd1 _14165_/X
+ sky130_fd_sc_hd__o211a_1
X_11377_ hold5735/X _11765_/B _11376_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11377_/X
+ sky130_fd_sc_hd__o211a_1
X_13116_ hold5294/X _13115_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__mux2_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ hold2056/X _16600_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__mux2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _15549_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13056_/C _13044_/X _13046_/X _09339_/A vssd1 vssd1 vccd1 vccd1 _13047_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _18053_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_1
X_10259_ hold2803/X hold4033/X _10643_/C vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__mux2_1
X_17855_ _17855_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
X_16806_ _18009_/CLK _16806_/D vssd1 vssd1 vccd1 vccd1 _16806_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_18__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_18__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_17786_ _17882_/CLK hold905/X vssd1 vssd1 vccd1 vccd1 hold904/A sky130_fd_sc_hd__dfxtp_1
X_14998_ _15213_/A _15018_/B vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__or2_1
X_16737_ _18069_/CLK _16737_/D vssd1 vssd1 vccd1 vccd1 _16737_/Q sky130_fd_sc_hd__dfxtp_1
X_13949_ hold2670/X _13980_/B _13948_/X _14147_/C1 vssd1 vssd1 vccd1 vccd1 _13949_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16668_ _18226_/CLK _16668_/D vssd1 vssd1 vccd1 vccd1 _16668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18407_ _18407_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15619_ _17282_/CLK _15619_/D vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _18221_/CLK _16599_/D vssd1 vssd1 vccd1 vccd1 _16599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ hold949/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__or2_1
X_18338_ _18397_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09071_ hold1140/X _09119_/A2 _09070_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _09071_/X
+ sky130_fd_sc_hd__o211a_1
X_18269_ _18339_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_272_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17901_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08022_ hold1606/X _08029_/B _08021_/X _08159_/A vssd1 vssd1 vccd1 vccd1 _08022_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 hold701/A vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 hold712/A vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_201_wb_clk_i clkbuf_5_19__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18033_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 hold789/X vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 hold750/X vssd1 vssd1 vccd1 vccd1 hold751/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold756 hold756/A vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold767 hold767/A vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 hold778/A vssd1 vssd1 vccd1 vccd1 input51/A sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ hold5118/X _10067_/B _09972_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
Xhold789 input42/X vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ hold44/X hold169/X _08932_/S vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__mux2_1
Xhold2102 _15577_/Q vssd1 vssd1 vccd1 vccd1 hold2102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2113 _15610_/Q vssd1 vssd1 vccd1 vccd1 hold2113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2124 _09320_/X vssd1 vssd1 vccd1 vccd1 _16270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 _18345_/Q vssd1 vssd1 vccd1 vccd1 hold2135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 _18386_/Q vssd1 vssd1 vccd1 vccd1 hold1401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2146 _08046_/X vssd1 vssd1 vccd1 vccd1 _15664_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _15473_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _16046_/D sky130_fd_sc_hd__and2_1
Xhold1412 _17965_/Q vssd1 vssd1 vccd1 vccd1 hold1412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2157 _18132_/Q vssd1 vssd1 vccd1 vccd1 hold2157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 _15601_/Q vssd1 vssd1 vccd1 vccd1 hold2168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 _07874_/X vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2179 _12645_/X vssd1 vssd1 vccd1 vccd1 _17391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _17857_/Q vssd1 vssd1 vccd1 vccd1 hold1434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1445 _15869_/Q vssd1 vssd1 vccd1 vccd1 hold1445/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1456 _08093_/X vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07806_ hold1504/X _07801_/B _09339_/B vssd1 vssd1 vccd1 vccd1 _07806_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08786_ _15473_/A hold97/X vssd1 vssd1 vccd1 vccd1 _16013_/D sky130_fd_sc_hd__and2_1
Xhold1467 _17512_/Q vssd1 vssd1 vccd1 vccd1 hold1467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 _18192_/Q vssd1 vssd1 vccd1 vccd1 hold1478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _18186_/Q vssd1 vssd1 vccd1 vccd1 hold1489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ _07804_/A _09447_/C _15334_/A _09406_/X vssd1 vssd1 vccd1 vccd1 _09407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09338_ hold2151/X _09338_/A2 _09337_/X _12927_/A vssd1 vssd1 vccd1 vccd1 _09338_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ hold335/X _16246_/Q _09277_/S vssd1 vssd1 vccd1 vccd1 hold336/A sky130_fd_sc_hd__mux2_1
X_11300_ _17772_/Q hold3799/X _12323_/C vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12280_ _12374_/A _12374_/B _12279_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ hold1034/X _16901_/Q _12305_/C vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ _16878_/Q _11201_/B _11201_/C vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__and3_1
Xhold4060 _09835_/X vssd1 vssd1 vccd1 vccd1 _16435_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10113_ _10563_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__or2_1
Xhold4071 _16673_/Q vssd1 vssd1 vccd1 vccd1 hold4071/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4082 _09574_/X vssd1 vssd1 vccd1 vccd1 _16348_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15970_ _17292_/CLK _15970_/D vssd1 vssd1 vccd1 vccd1 hold392/A sky130_fd_sc_hd__dfxtp_1
Xhold4093 _16553_/Q vssd1 vssd1 vccd1 vccd1 hold4093/X sky130_fd_sc_hd__dlygate4sd3_1
X_11093_ hold2580/X _16855_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3370 _17151_/Q vssd1 vssd1 vccd1 vccd1 hold3370/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ _13230_/A _10098_/A _10043_/X vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__a21oi_1
X_14921_ hold2923/X _14952_/B _14920_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _14921_/X
+ sky130_fd_sc_hd__o211a_1
Xhold3381 _12947_/X vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3392 _16964_/Q vssd1 vssd1 vccd1 vccd1 hold3392/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_leaf_77_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17523_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__buf_4
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2680 _18296_/Q vssd1 vssd1 vccd1 vccd1 hold2680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _17738_/CLK _17640_/D vssd1 vssd1 vccd1 vccd1 _17640_/Q sky130_fd_sc_hd__dfxtp_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _15191_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__or2_1
Xhold2691 _18083_/Q vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1990 _15749_/Q vssd1 vssd1 vccd1 vccd1 hold1990/X sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ hold3907/X _13710_/A _13802_/X vssd1 vssd1 vccd1 vccd1 _13803_/Y sky130_fd_sc_hd__a21oi_1
X_14783_ hold2322/X _14774_/B _14782_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14783_/X
+ sky130_fd_sc_hd__o211a_1
X_17571_ _17731_/CLK _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
X_11995_ hold4553/X _12377_/B _11994_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _11995_/X
+ sky130_fd_sc_hd__o211a_1
X_13734_ _13734_/A _13734_/B vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__or2_1
X_16522_ _18176_/CLK _16522_/D vssd1 vssd1 vccd1 vccd1 _16522_/Q sky130_fd_sc_hd__dfxtp_1
X_10946_ hold1778/X _16806_/Q _11717_/C vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16453_ _18373_/CLK _16453_/D vssd1 vssd1 vccd1 vccd1 _16453_/Q sky130_fd_sc_hd__dfxtp_1
X_13665_ _13776_/A _13665_/B vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__or2_1
X_10877_ hold399/X hold5679/X _11201_/C vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_128_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15482_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__and2_1
X_12616_ hold995/X hold3020/X _12676_/S vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__mux2_1
X_16384_ _18330_/CLK _16384_/D vssd1 vssd1 vccd1 vccd1 _16384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13788_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__or2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18123_ _18233_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
X_15335_ hold687/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ hold1172/X _17360_/Q _12922_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _17330_/Q _09362_/C _09362_/D hold691/X vssd1 vssd1 vccd1 vccd1 _15266_/X
+ sky130_fd_sc_hd__a22o_1
X_18054_ _18054_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12478_ _17332_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _13308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17005_ _17856_/CLK _17005_/D vssd1 vssd1 vccd1 vccd1 _17005_/Q sky130_fd_sc_hd__dfxtp_1
X_14217_ _14897_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__or2_2
X_11429_ hold2620/X _16967_/Q _12299_/C vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__mux2_1
X_15197_ _15197_/A _15211_/B vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _15547_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14079_ hold1265/X _14094_/B _14078_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _14079_/X
+ sky130_fd_sc_hd__o211a_1
X_17907_ _17907_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_1
X_08640_ _12428_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _15942_/D sky130_fd_sc_hd__and2_1
X_17838_ _17870_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _12428_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _15909_/D sky130_fd_sc_hd__and2_1
X_17769_ _17769_/CLK hold737/X vssd1 vssd1 vccd1 vccd1 _17769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _07788_/A _09120_/Y hold802/X _18459_/Q vssd1 vssd1 vccd1 vccd1 hold803/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09054_ hold44/X hold462/X _09056_/S vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_142_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08005_ _15519_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 hold531/A vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold553 hold553/A vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 hold564/A vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold575 hold575/A vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 hold586/A vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold597/A vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09956_ hold1317/X _16476_/Q _10271_/S vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__mux2_1
X_08907_ _12422_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _16071_/D sky130_fd_sc_hd__and2_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ hold2478/X hold5352/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__mux2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _18253_/Q vssd1 vssd1 vccd1 vccd1 hold1220/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _15620_/Q vssd1 vssd1 vccd1 vccd1 hold1231/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ hold184/X hold718/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__mux2_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _15776_/Q vssd1 vssd1 vccd1 vccd1 hold1242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _17841_/Q vssd1 vssd1 vccd1 vccd1 hold1253/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 _09135_/X vssd1 vssd1 vccd1 vccd1 _16180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 _15780_/Q vssd1 vssd1 vccd1 vccd1 hold1275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _18356_/Q vssd1 vssd1 vccd1 vccd1 hold1286/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ hold17/X _16005_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 hold1297/A vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _10998_/A _10800_/B vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _17084_/Q _12323_/B _12323_/C vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__and3_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _11667_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_194_wb_clk_i clkbuf_5_24__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13450_ hold4437/X _13832_/B _13449_/X _08379_/A vssd1 vssd1 vccd1 vccd1 _13450_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10662_ _11061_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__or2_1
X_12401_ hold53/X hold186/X _12439_/S vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_wb_clk_i clkbuf_5_25__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18267_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ hold5168/X _13859_/B _13380_/X _08387_/A vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ _16528_/Q _10521_/A _10592_/X vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__a21oi_1
X_15120_ hold2372/X _15113_/B _15119_/X _15066_/A vssd1 vssd1 vccd1 vccd1 _15120_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12332_ _17268_/Q _12362_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15105_/A hold980/X _15069_/S vssd1 vssd1 vccd1 vccd1 hold981/A sky130_fd_sc_hd__mux2_1
X_12263_ hold2102/X _17245_/Q _13388_/S vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__mux2_1
X_14002_ hold944/X _14052_/B vssd1 vssd1 vccd1 vccd1 _14002_/X sky130_fd_sc_hd__or2_1
X_11214_ hold5266/X _11103_/A _11213_/X vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__a21oi_1
X_12194_ hold1792/X hold4261/X _13796_/S vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput73 _13137_/A vssd1 vssd1 vccd1 vccd1 output73/X sky130_fd_sc_hd__buf_6
X_11145_ hold3751/X _11637_/A _11144_/X vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__a21oi_1
Xoutput84 _13217_/A vssd1 vssd1 vccd1 vccd1 output84/X sky130_fd_sc_hd__buf_6
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput95 _13297_/A vssd1 vssd1 vccd1 vccd1 output95/X sky130_fd_sc_hd__buf_6
X_15953_ _17300_/CLK _15953_/D vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__dfxtp_1
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__or2_1
X_10027_ _11203_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__nor2_1
X_14904_ hold667/A _14910_/B vssd1 vssd1 vccd1 vccd1 hold638/A sky130_fd_sc_hd__or2_1
X_15884_ _17723_/CLK _15884_/D vssd1 vssd1 vccd1 vccd1 _15884_/Q sky130_fd_sc_hd__dfxtp_1
X_17623_ _17719_/CLK _17623_/D vssd1 vssd1 vccd1 vccd1 _17623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ hold2584/X _14828_/B _14834_/X _15003_/C1 vssd1 vssd1 vccd1 vccd1 _14835_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _18229_/CLK _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14766_ _15213_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__or2_1
X_11978_ hold2207/X hold4423/X _13871_/C vssd1 vssd1 vccd1 vccd1 _11979_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_187_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16505_ _18358_/CLK _16505_/D vssd1 vssd1 vccd1 vccd1 _16505_/Q sky130_fd_sc_hd__dfxtp_1
X_13717_ hold4995/X _13811_/B _13716_/X _15534_/C1 vssd1 vssd1 vccd1 vccd1 _13717_/X
+ sky130_fd_sc_hd__o211a_1
X_10929_ _11121_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__or2_1
X_17485_ _17485_/CLK _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/Q sky130_fd_sc_hd__dfxtp_1
X_14697_ hold1673/X _14720_/B _14696_/X _14833_/C1 vssd1 vssd1 vccd1 vccd1 _14697_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16436_ _18381_/CLK _16436_/D vssd1 vssd1 vccd1 vccd1 _16436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ hold4526/X _13856_/B _13647_/X _08381_/A vssd1 vssd1 vccd1 vccd1 _13648_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _18416_/CLK _16367_/D vssd1 vssd1 vccd1 vccd1 _16367_/Q sky130_fd_sc_hd__dfxtp_1
X_13579_ hold3344/X _13823_/B _13578_/X _13771_/C1 vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18106_ _18140_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15318_ hold382/X _15484_/A2 _15451_/A2 hold457/X vssd1 vssd1 vccd1 vccd1 _15318_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _16314_/CLK _16298_/D vssd1 vssd1 vccd1 vccd1 _16298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5508 _16809_/Q vssd1 vssd1 vccd1 vccd1 hold5508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5519 _10834_/X vssd1 vssd1 vccd1 vccd1 _16768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ _18069_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15249_ hold549/X _15485_/A2 _15447_/B1 hold446/X _15248_/X vssd1 vssd1 vccd1 vccd1
+ _15252_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4807 _17722_/Q vssd1 vssd1 vccd1 vccd1 hold4807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4818 _17175_/Q vssd1 vssd1 vccd1 vccd1 hold4818/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4829 _13333_/X vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09810_ _09948_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout307 fanout337/X vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__clkbuf_4
Xfanout318 _10998_/A vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__buf_4
Xfanout329 _10098_/A vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__clkbuf_4
X_09741_ _09933_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__or2_1
X_09672_ _09954_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__or2_1
XFILLER_0_154_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08623_ hold81/X hold726/X _08661_/S vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ hold136/X hold339/X _08594_/S vssd1 vssd1 vccd1 vccd1 hold340/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ hold2153/X _08488_/B _08484_/Y _08379_/A vssd1 vssd1 vccd1 vccd1 _08485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09106_ _15221_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09037_ _15374_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _16135_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 hold361/A vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold394/A vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout830 _14859_/C1 vssd1 vssd1 vccd1 vccd1 _14849_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout841 fanout842/X vssd1 vssd1 vccd1 vccd1 fanout841/X sky130_fd_sc_hd__buf_4
Xfanout852 _11791_/A vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__buf_6
X_09939_ _09987_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__or2_1
Xfanout863 _15215_/A vssd1 vssd1 vccd1 vccd1 _15000_/A sky130_fd_sc_hd__buf_12
Xfanout874 hold616/X vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__buf_4
Xfanout885 _15195_/A vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__buf_6
Xfanout896 _14850_/A vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__buf_8
XFILLER_0_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12950_ hold3596/X _12949_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__mux2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _08073_/X vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _12018_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__or2_1
Xhold1061 _17949_/Q vssd1 vssd1 vccd1 vccd1 hold1061/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 _13942_/X vssd1 vssd1 vccd1 vccd1 _13943_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 _14071_/X vssd1 vssd1 vccd1 vccd1 _17840_/D sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ hold3246/X _12880_/X _12920_/S vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _15562_/Q vssd1 vssd1 vccd1 vccd1 hold1094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14728_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14620_/X sky130_fd_sc_hd__or2_1
X_11832_ _13794_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__or2_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_304_wb_clk_i clkbuf_5_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14551_ _15231_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14551_/X sky130_fd_sc_hd__or2_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ hold5324/X _11694_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13502_ hold977/X _17621_/Q _13886_/C vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ hold5596/X _10897_/A2 _10713_/X _14813_/C1 vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__o211a_1
X_17270_ _17906_/CLK _17270_/D vssd1 vssd1 vccd1 vccd1 _17270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ hold2068/X _14481_/B _14481_/Y _14548_/C1 vssd1 vssd1 vccd1 vccd1 _14482_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ _11694_/A _11694_/B vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__or2_1
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13433_ hold1187/X hold3293/X _13862_/C vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__mux2_1
X_16221_ _17453_/CLK _16221_/D vssd1 vssd1 vccd1 vccd1 _16221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _11218_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16152_ _17517_/CLK _16152_/D vssd1 vssd1 vccd1 vccd1 _16152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13364_ hold908/X hold3902/X _13844_/C vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10576_ _11194_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _10576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15103_ _15103_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__or2_1
XFILLER_0_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12315_ hold3773/X _12285_/A _12314_/X vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16083_ _17751_/CLK _16083_/D vssd1 vssd1 vccd1 vccd1 hold532/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _13311_/A1 _13293_/X _13294_/X _13311_/C1 vssd1 vssd1 vccd1 vccd1 _13295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15052_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15034_/X sky130_fd_sc_hd__and2_1
X_12246_ _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_91_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17302_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ _12279_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_5_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17475_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11128_ hold5674/X _11789_/B _11127_/X _14350_/A vssd1 vssd1 vccd1 vccd1 _11128_/X
+ sky130_fd_sc_hd__o211a_1
X_16985_ _17769_/CLK _16985_/D vssd1 vssd1 vccd1 vccd1 _16985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15936_ _18425_/CLK _15936_/D vssd1 vssd1 vccd1 vccd1 hold543/A sky130_fd_sc_hd__dfxtp_1
X_11059_ hold5606/X _11156_/B _11058_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _11059_/X
+ sky130_fd_sc_hd__o211a_1
X_15867_ _17738_/CLK _15867_/D vssd1 vssd1 vccd1 vccd1 _15867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ _17734_/CLK _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14818_ _15103_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__or2_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _17697_/CLK _15798_/D vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _18380_/CLK _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14749_ hold2911/X _14772_/B _14748_/X _14869_/C1 vssd1 vssd1 vccd1 vccd1 _14749_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _15549_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17482_/CLK _17468_/D vssd1 vssd1 vccd1 vccd1 _17468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16419_ _18388_/CLK _16419_/D vssd1 vssd1 vccd1 vccd1 _16419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17399_ _18451_/CLK _17399_/D vssd1 vssd1 vccd1 vccd1 _17399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6006 la_data_in[1] vssd1 vssd1 vccd1 vccd1 hold888/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold6017 _16307_/Q vssd1 vssd1 vccd1 vccd1 hold6017/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6028 _16309_/Q vssd1 vssd1 vccd1 vccd1 hold6028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6039 data_in[10] vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold5305 _10024_/Y vssd1 vssd1 vccd1 vccd1 _16498_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5316 _10017_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5327 _16367_/Q vssd1 vssd1 vccd1 vccd1 hold5327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5338 _16364_/Q vssd1 vssd1 vccd1 vccd1 hold5338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5349 _11851_/X vssd1 vssd1 vccd1 vccd1 _17107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4604 _11254_/X vssd1 vssd1 vccd1 vccd1 _16908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4615 _17035_/Q vssd1 vssd1 vccd1 vccd1 hold4615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4626 _10729_/X vssd1 vssd1 vccd1 vccd1 _16733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4637 _17157_/Q vssd1 vssd1 vccd1 vccd1 hold4637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3903 _13845_/Y vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold4648 _11512_/X vssd1 vssd1 vccd1 vccd1 _16994_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3914 _10567_/Y vssd1 vssd1 vccd1 vccd1 _16679_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4659 _16872_/Q vssd1 vssd1 vccd1 vccd1 hold4659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3925 _10426_/X vssd1 vssd1 vccd1 vccd1 _16632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3936 _16632_/Q vssd1 vssd1 vccd1 vccd1 hold3936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3947 _13873_/Y vssd1 vssd1 vccd1 vccd1 _17744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3958 _09949_/X vssd1 vssd1 vccd1 vccd1 _16473_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3969 _17587_/Q vssd1 vssd1 vccd1 vccd1 hold3969/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout148 _12800_/S vssd1 vssd1 vccd1 vccd1 _12806_/S sky130_fd_sc_hd__clkbuf_8
Xfanout159 _13808_/B vssd1 vssd1 vccd1 vccd1 _13805_/B sky130_fd_sc_hd__buf_4
X_07985_ hold2392/X _07978_/B _07984_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _07985_/X
+ sky130_fd_sc_hd__o211a_1
X_09724_ hold3888/X _10028_/B _09723_/X _15052_/A vssd1 vssd1 vccd1 vccd1 _09724_/X
+ sky130_fd_sc_hd__o211a_1
X_09655_ hold4528/X _10049_/B _09654_/X _14939_/C1 vssd1 vssd1 vccd1 vccd1 _09655_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08606_ _08970_/A _08606_/B vssd1 vssd1 vccd1 vccd1 _15925_/D sky130_fd_sc_hd__and2_1
XFILLER_0_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09586_ hold5171/X _10628_/B _09585_/X _15024_/A vssd1 vssd1 vccd1 vccd1 _09586_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08537_ _15354_/A hold641/X vssd1 vssd1 vccd1 vccd1 _15892_/D sky130_fd_sc_hd__and2_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ hold883/X _08500_/B vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08399_ _15513_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ hold1478/X _16634_/Q _10649_/C vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ hold2300/X hold3247/X _10640_/C vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12100_ hold4261/X _12308_/B _12099_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _12100_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13080_ _13073_/X _13079_/X _13048_/A vssd1 vssd1 vccd1 vccd1 _17528_/D sky130_fd_sc_hd__o21a_1
Xhold5850 _16282_/Q vssd1 vssd1 vccd1 vccd1 hold5850/X sky130_fd_sc_hd__dlygate4sd3_1
X_10292_ hold1615/X hold4143/X _10625_/C vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__mux2_1
Xhold5861 hold5861/A vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_12
Xhold5872 _18425_/Q vssd1 vssd1 vccd1 vccd1 hold5872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5883 _16175_/Q vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__buf_1
X_12031_ hold4899/X _12356_/B _12030_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12031_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5894 _16320_/Q vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout660 fanout842/X vssd1 vssd1 vccd1 vccd1 fanout660/X sky130_fd_sc_hd__buf_4
XFILLER_0_176_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout671 _08137_/A vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__buf_2
XFILLER_0_189_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout682 _14171_/C1 vssd1 vssd1 vccd1 vccd1 _14193_/C1 sky130_fd_sc_hd__buf_4
X_16770_ _18032_/CLK _16770_/D vssd1 vssd1 vccd1 vccd1 _16770_/Q sky130_fd_sc_hd__dfxtp_1
X_13982_ _15109_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13982_/Y sky130_fd_sc_hd__nand2_1
Xfanout693 _15244_/A vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__clkbuf_4
X_15721_ _17128_/CLK _15721_/D vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12933_ _12933_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _17487_/D sky130_fd_sc_hd__and2_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _18454_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _17260_/CLK _15652_/D vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12924_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _17464_/D sky130_fd_sc_hd__and2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ hold1844/X _14610_/B _14602_/X _14955_/C1 vssd1 vssd1 vccd1 vccd1 _14603_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ hold3249/X _12302_/B _11814_/X _12831_/A vssd1 vssd1 vccd1 vccd1 _11815_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18371_/CLK hold959/X vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15583_ _17283_/CLK _15583_/D vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfxtp_1
X_12795_ _12825_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _17441_/D sky130_fd_sc_hd__and2_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17531_/CLK hold27/X vssd1 vssd1 vccd1 vccd1 _17322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _12301_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11746_/Y sky130_fd_sc_hd__nor2_1
X_14534_ hold1244/X _14554_/A2 _14533_/X _13911_/A vssd1 vssd1 vccd1 vccd1 _14534_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _17253_/CLK _17253_/D vssd1 vssd1 vccd1 vccd1 _17253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11677_ hold5395/X _12338_/B _11676_/X _13923_/A vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__o211a_1
X_14465_ _14984_/A _14499_/B vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _17435_/CLK _16204_/D vssd1 vssd1 vccd1 vccd1 _16204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ _16700_/Q _10628_/B _10628_/C vssd1 vssd1 vccd1 vccd1 _10628_/X sky130_fd_sc_hd__and3_1
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13416_ _13800_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13416_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17184_ _17216_/CLK _17184_/D vssd1 vssd1 vccd1 vccd1 _17184_/Q sky130_fd_sc_hd__dfxtp_1
X_14396_ hold2913/X hold209/X _14395_/X _14384_/A vssd1 vssd1 vccd1 vccd1 _14396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16135_ _17287_/CLK _16135_/D vssd1 vssd1 vccd1 vccd1 hold724/A sky130_fd_sc_hd__dfxtp_1
X_13347_ _13737_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__or2_1
X_10559_ hold1702/X _16677_/Q _10568_/C vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ _13278_/A _13310_/B vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__or2_1
X_16066_ _18408_/CLK _16066_/D vssd1 vssd1 vccd1 vccd1 hold563/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15017_ hold1368/X _15004_/B _15016_/X _15216_/C1 vssd1 vssd1 vccd1 vccd1 _15017_/X
+ sky130_fd_sc_hd__o211a_1
X_12229_ hold4677/X _12323_/B _12228_/X _13929_/A vssd1 vssd1 vccd1 vccd1 _12229_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2509 _17845_/Q vssd1 vssd1 vccd1 vccd1 hold2509/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1808 _08269_/X vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 _14145_/X vssd1 vssd1 vccd1 vccd1 _17876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_297_wb_clk_i clkbuf_5_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17686_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16968_ _17880_/CLK _16968_/D vssd1 vssd1 vccd1 vccd1 _16968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_226_wb_clk_i clkbuf_5_22__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17905_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15919_ _18410_/CLK _15919_/D vssd1 vssd1 vccd1 vccd1 hold645/A sky130_fd_sc_hd__dfxtp_1
X_16899_ _18070_/CLK _16899_/D vssd1 vssd1 vccd1 vccd1 _16899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09440_ _18463_/A _15314_/A vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__and2_1
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ hold348/X _09362_/C _09386_/D hold651/X _09370_/X vssd1 vssd1 vccd1 vccd1
+ _09375_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08322_ hold1822/X _08323_/B _08321_/Y _13801_/C1 vssd1 vssd1 vccd1 vccd1 _08322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08253_ hold1177/X _08262_/B _08252_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _08253_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ hold985/X _08209_/B _08183_/X _08371_/A vssd1 vssd1 vccd1 vccd1 hold986/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5102 _17715_/Q vssd1 vssd1 vccd1 vccd1 hold5102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5113 _11977_/X vssd1 vssd1 vccd1 vccd1 _17149_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5124 _17683_/Q vssd1 vssd1 vccd1 vccd1 hold5124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold5135 _09595_/X vssd1 vssd1 vccd1 vccd1 _16355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5146 _17649_/Q vssd1 vssd1 vccd1 vccd1 hold5146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4401 _17067_/Q vssd1 vssd1 vccd1 vccd1 hold4401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4412 _13723_/X vssd1 vssd1 vccd1 vccd1 _17694_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold5157 _13669_/X vssd1 vssd1 vccd1 vccd1 _17676_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5168 _17612_/Q vssd1 vssd1 vccd1 vccd1 hold5168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4423 _17150_/Q vssd1 vssd1 vccd1 vccd1 hold4423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4434 _12208_/X vssd1 vssd1 vccd1 vccd1 _17226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3700 _10647_/Y vssd1 vssd1 vccd1 vccd1 _10648_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold5179 _17642_/Q vssd1 vssd1 vccd1 vccd1 hold5179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4445 _17182_/Q vssd1 vssd1 vccd1 vccd1 hold4445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3711 _16462_/Q vssd1 vssd1 vccd1 vccd1 hold3711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4456 _11245_/X vssd1 vssd1 vccd1 vccd1 _16905_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3722 _16345_/Q vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold4467 _16413_/Q vssd1 vssd1 vccd1 vccd1 hold4467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3733 _12364_/Y vssd1 vssd1 vccd1 vccd1 _17278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4478 _11701_/X vssd1 vssd1 vccd1 vccd1 _17057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3744 _11737_/Y vssd1 vssd1 vccd1 vccd1 _17069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4489 _10873_/X vssd1 vssd1 vccd1 vccd1 _16781_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3755 _10621_/Y vssd1 vssd1 vccd1 vccd1 _16697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3766 _13819_/Y vssd1 vssd1 vccd1 vccd1 _17726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3777 _12298_/Y vssd1 vssd1 vccd1 vccd1 _17256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3788 _11724_/Y vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold3799 _16924_/Q vssd1 vssd1 vccd1 vccd1 hold3799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07968_ _15537_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__or2_1
X_09707_ hold2262/X hold5516/X _09998_/C vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ hold2674/X _07918_/B _07898_/X _08135_/A vssd1 vssd1 vccd1 vccd1 _07899_/X
+ sky130_fd_sc_hd__o211a_1
X_09638_ hold1698/X hold5639/X _10022_/C vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09569_ hold1430/X _13246_/A _10271_/S vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ hold1734/X hold4277/X _11792_/C vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ hold1459/X hold2925/X _12982_/S vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ hold1998/X hold4367/X _11726_/C vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_191_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14250_ _14984_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__or2_1
X_11462_ hold2241/X hold5435/X _11753_/C vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ _13201_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10413_ _10551_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10413_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ hold1204/X _14202_/B _14180_/X _14203_/C1 vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__o211a_1
X_11393_ hold2193/X _16955_/Q _12323_/C vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__mux2_1
X_13132_ hold3665/X _13131_/X _13244_/S vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_2
X_10344_ _10542_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__or2_1
XFILLER_0_143_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ _18069_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_1
Xhold5680 _10783_/X vssd1 vssd1 vccd1 vccd1 _16751_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13063_ _13183_/A1 _13061_/X _13062_/X _13183_/C1 vssd1 vssd1 vccd1 vccd1 _13063_/X
+ sky130_fd_sc_hd__o211a_1
Xhold5691 _16854_/Q vssd1 vssd1 vccd1 vccd1 hold5691/X sky130_fd_sc_hd__dlygate4sd3_1
X_10275_ _10563_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__or2_1
X_12014_ hold1105/X hold4218/X _13811_/C vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__mux2_1
Xhold4990 _17213_/Q vssd1 vssd1 vccd1 vccd1 hold4990/X sky130_fd_sc_hd__dlygate4sd3_1
X_17871_ _17903_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _18025_/CLK _16822_/D vssd1 vssd1 vccd1 vccd1 _16822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout490 _10874_/S vssd1 vssd1 vccd1 vccd1 _10022_/C sky130_fd_sc_hd__clkbuf_8
Xclkbuf_5_17__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_5_17__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_16753_ _18053_/CLK _16753_/D vssd1 vssd1 vccd1 vccd1 _16753_/Q sky130_fd_sc_hd__dfxtp_1
X_13965_ hold2597/X _13980_/B _13964_/X _14510_/C1 vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _17282_/CLK _15704_/D vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ hold2590/X _17483_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16684_ _18210_/CLK _16684_/D vssd1 vssd1 vccd1 vccd1 _16684_/Q sky130_fd_sc_hd__dfxtp_1
X_13896_ hold892/X hold1088/X hold244/X vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__mux2_1
X_18423_ _18423_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ _17211_/CLK _15635_/D vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ hold2530/X _17460_/Q _12919_/S vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__mux2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18378_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15566_ _17902_/CLK _15566_/D vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ hold1599/X _17437_/Q _12820_/S vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _18421_/CLK _17305_/D vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _14517_/A _14545_/B vssd1 vssd1 vccd1 vccd1 _14517_/X sky130_fd_sc_hd__or2_1
XFILLER_0_185_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18285_ _18363_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _17067_/Q _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__and3_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15497_ _14972_/A hold1780/X _15505_/S vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_153_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _17268_/CLK _17236_/D vssd1 vssd1 vccd1 vccd1 _17236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448_ hold607/X hold273/A vssd1 vssd1 vccd1 vccd1 _14479_/B sky130_fd_sc_hd__or2_4
XFILLER_0_126_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17167_ _17263_/CLK _17167_/D vssd1 vssd1 vccd1 vccd1 _17167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 hold905/A vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ hold173/X hold422/X hold275/X vssd1 vssd1 vccd1 vccd1 hold423/A sky130_fd_sc_hd__mux2_1
Xhold916 hold916/A vssd1 vssd1 vccd1 vccd1 hold916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 hold927/A vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__clkbuf_2
X_16118_ _17341_/CLK _16118_/D vssd1 vssd1 vccd1 vccd1 hold646/A sky130_fd_sc_hd__dfxtp_1
Xhold938 hold938/A vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17098_ _18445_/CLK _17098_/D vssd1 vssd1 vccd1 vccd1 _17098_/Q sky130_fd_sc_hd__dfxtp_1
Xhold949 hold949/A vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__buf_8
Xhold3007 _12911_/X vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__dlygate4sd3_1
X_16049_ _17525_/CLK _16049_/D vssd1 vssd1 vccd1 vccd1 hold695/A sky130_fd_sc_hd__dfxtp_1
X_08940_ _12442_/A hold613/X vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3018 _17474_/Q vssd1 vssd1 vccd1 vccd1 hold3018/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3029 _18138_/Q vssd1 vssd1 vccd1 vccd1 hold3029/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2306 _18150_/Q vssd1 vssd1 vccd1 vccd1 hold2306/X sky130_fd_sc_hd__dlygate4sd3_1
X_08871_ _12428_/A hold286/X vssd1 vssd1 vccd1 vccd1 _16053_/D sky130_fd_sc_hd__and2_1
Xhold2317 _07931_/X vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2328 _17804_/Q vssd1 vssd1 vccd1 vccd1 hold2328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 _14424_/X vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 _08218_/X vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07822_ hold173/X hold335/X vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__or2_1
Xhold1616 _14709_/X vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 _17880_/Q vssd1 vssd1 vccd1 vccd1 hold1627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 _15779_/Q vssd1 vssd1 vccd1 vccd1 hold1638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 _09310_/X vssd1 vssd1 vccd1 vccd1 _16265_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09423_ _07804_/A _09463_/A _15334_/A _09422_/X vssd1 vssd1 vccd1 vccd1 _09423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _09400_/A _09366_/B _09361_/C vssd1 vssd1 vccd1 vccd1 _09354_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_164_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ hold747/X _08305_/B vssd1 vssd1 vccd1 vccd1 _08305_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09285_ _14913_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _14850_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__or2_1
XFILLER_0_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ _08355_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _15557_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__or2_1
Xhold4220 _17603_/Q vssd1 vssd1 vccd1 vccd1 hold4220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4231 _13537_/X vssd1 vssd1 vccd1 vccd1 _17632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4242 _16602_/Q vssd1 vssd1 vccd1 vccd1 hold4242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4253 _10495_/X vssd1 vssd1 vccd1 vccd1 _16655_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4264 _10516_/X vssd1 vssd1 vccd1 vccd1 _16662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3530 _09967_/X vssd1 vssd1 vccd1 vccd1 _16479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_148_wb_clk_i clkbuf_5_30__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18095_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold4275 _16440_/Q vssd1 vssd1 vccd1 vccd1 hold4275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4286 _10336_/X vssd1 vssd1 vccd1 vccd1 _16602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3541 _17431_/Q vssd1 vssd1 vccd1 vccd1 hold3541/X sky130_fd_sc_hd__dlygate4sd3_1
X_10060_ _11194_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__nor2_1
Xhold3552 _17647_/Q vssd1 vssd1 vccd1 vccd1 hold3552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4297 _16612_/Q vssd1 vssd1 vccd1 vccd1 hold4297/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3563 _09559_/X vssd1 vssd1 vccd1 vccd1 _16343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3574 _13588_/X vssd1 vssd1 vccd1 vccd1 _17649_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2840 _15691_/Q vssd1 vssd1 vccd1 vccd1 hold2840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3585 _12929_/X vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2851 _16161_/Q vssd1 vssd1 vccd1 vccd1 hold2851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3596 _17493_/Q vssd1 vssd1 vccd1 vccd1 hold3596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2862 _18056_/Q vssd1 vssd1 vccd1 vccd1 hold2862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2873 _14587_/X vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2884 _18092_/Q vssd1 vssd1 vccd1 vccd1 hold2884/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2895 _17783_/Q vssd1 vssd1 vccd1 vccd1 hold2895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13750_ hold4708/X _13844_/B _13749_/X _08151_/A vssd1 vssd1 vccd1 vccd1 _13750_/X
+ sky130_fd_sc_hd__o211a_1
X_10962_ _11136_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10962_/X sky130_fd_sc_hd__or2_1
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ hold3410/X _12700_/X _12821_/S vssd1 vssd1 vccd1 vccd1 _12701_/X sky130_fd_sc_hd__mux2_1
X_13681_ hold4731/X _13868_/B _13680_/X _13681_/C1 vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__o211a_1
X_10893_ _11097_/A _10893_/B vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__or2_1
XFILLER_0_168_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15420_ hold527/X _09365_/B _15485_/B1 hold388/X _15418_/X vssd1 vssd1 vccd1 vccd1
+ _15422_/C sky130_fd_sc_hd__a221o_1
X_12632_ hold3072/X _12631_/X _12677_/S vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_182_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15351_ _16299_/Q _09362_/A _09392_/B hold612/X _15350_/X vssd1 vssd1 vccd1 vccd1
+ _15352_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12563_ hold3588/X _12562_/X _12953_/S vssd1 vssd1 vccd1 vccd1 _12563_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _12246_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__or2_1
X_14302_ hold949/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14302_/X sky130_fd_sc_hd__or2_1
X_18070_ _18070_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
X_15282_ _15489_/A _15282_/B _15282_/C _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/X
+ sky130_fd_sc_hd__or4_1
X_12494_ _17340_/Q _12508_/B vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17021_ _17891_/CLK _17021_/D vssd1 vssd1 vccd1 vccd1 _17021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11616_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__or2_1
X_14233_ _14913_/A hold273/A vssd1 vssd1 vccd1 vccd1 _14280_/B sky130_fd_sc_hd__or2_4
XFILLER_0_150_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14164_ _14218_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__or2_1
X_11376_ _11670_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ hold3261/X _10637_/B _10326_/X _14877_/C1 vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o211a_1
X_13115_ _13114_/X hold3737/X _13251_/S vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__mux2_1
X_14095_ hold2066/X _14094_/B _14094_/Y _13897_/A vssd1 vssd1 vccd1 vccd1 _14095_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _13053_/A _13046_/C _13046_/D vssd1 vssd1 vccd1 vccd1 _13046_/X
+ sky130_fd_sc_hd__or4_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17923_/CLK _17923_/D vssd1 vssd1 vccd1 vccd1 _17923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10258_ hold4365/X _10640_/B _10257_/X _14883_/C1 vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ _18051_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_1
X_10189_ hold4232/X _10465_/A2 _10188_/X _14941_/C1 vssd1 vssd1 vccd1 vccd1 _10189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ _18042_/CLK _16805_/D vssd1 vssd1 vccd1 vccd1 _16805_/Q sky130_fd_sc_hd__dfxtp_1
X_17785_ _17785_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
X_14997_ hold2234/X _15004_/B _14996_/X _15062_/A vssd1 vssd1 vccd1 vccd1 _14997_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16736_ _18035_/CLK _16736_/D vssd1 vssd1 vccd1 vccd1 _16736_/Q sky130_fd_sc_hd__dfxtp_1
X_13948_ _14218_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16667_ _18225_/CLK _16667_/D vssd1 vssd1 vccd1 vccd1 _16667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ _13888_/A _13879_/B vssd1 vssd1 vccd1 vccd1 _13879_/Y sky130_fd_sc_hd__nor2_1
X_18406_ _18406_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
X_15618_ _17584_/CLK _15618_/D vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfxtp_1
X_16598_ _18216_/CLK _16598_/D vssd1 vssd1 vccd1 vccd1 _16598_/Q sky130_fd_sc_hd__dfxtp_1
X_18337_ _18337_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15549_ _15549_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ hold892/X _09118_/B vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18268_ _18268_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _08311_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _17283_/CLK _17219_/D vssd1 vssd1 vccd1 vccd1 _17219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199_ _18231_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 hold724/A vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold735 hold735/A vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__buf_12
Xhold746 hold752/X vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 hold757/A vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 hold777/X vssd1 vssd1 vccd1 vccd1 hold778/A sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _10506_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__or2_1
Xhold779 input51/X vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_241_wb_clk_i clkbuf_5_20__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17715_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08923_ _15374_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _16079_/D sky130_fd_sc_hd__and2_1
Xhold2103 _07864_/X vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2114 _07933_/X vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2125 _17799_/Q vssd1 vssd1 vccd1 vccd1 hold2125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2136 _15122_/X vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1402 _15208_/X vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2147 _17821_/Q vssd1 vssd1 vccd1 vccd1 hold2147/X sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ hold50/X hold323/X _08860_/S vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1413 _14331_/X vssd1 vssd1 vccd1 vccd1 _17965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 _14679_/X vssd1 vssd1 vccd1 vccd1 _18132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 _18055_/Q vssd1 vssd1 vccd1 vccd1 hold1424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 _07915_/X vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 _14105_/X vssd1 vssd1 vccd1 vccd1 _17857_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07805_/Y sky130_fd_sc_hd__inv_2
Xhold1446 _08481_/X vssd1 vssd1 vccd1 vccd1 _15869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ hold44/X _16013_/Q _08793_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _15626_/Q vssd1 vssd1 vccd1 vccd1 hold1457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _13008_/X vssd1 vssd1 vccd1 vccd1 _17512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 _14805_/X vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09406_ _09438_/B _16289_/Q vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09337_ _15559_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _09272_/A hold236/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__and2_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08219_ _14726_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ hold2662/X _09218_/B _09198_/X _12813_/A vssd1 vssd1 vccd1 vccd1 _09199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ hold4875/X _12320_/B _11229_/X _13905_/A vssd1 vssd1 vccd1 vccd1 _11230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _12301_/A _11161_/B vssd1 vssd1 vccd1 vccd1 _11161_/Y sky130_fd_sc_hd__nor2_1
Xhold4050 _13609_/X vssd1 vssd1 vccd1 vccd1 _17656_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold4061 _16635_/Q vssd1 vssd1 vccd1 vccd1 hold4061/X sky130_fd_sc_hd__dlygate4sd3_1
X_10112_ hold2999/X _16528_/Q _10565_/C vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__mux2_1
Xhold4072 _10453_/X vssd1 vssd1 vccd1 vccd1 _16641_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11092_ hold5645/X _11213_/B _11091_/X _14879_/C1 vssd1 vssd1 vccd1 vccd1 _11092_/X
+ sky130_fd_sc_hd__o211a_1
Xhold4083 _16565_/Q vssd1 vssd1 vccd1 vccd1 hold4083/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold4094 _10093_/X vssd1 vssd1 vccd1 vccd1 _16521_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold3360 _16569_/Q vssd1 vssd1 vccd1 vccd1 hold3360/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ _16505_/Q _10601_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__and3_1
X_14920_ _15189_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__or2_1
Xhold3371 _11887_/X vssd1 vssd1 vccd1 vccd1 _17119_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3382 _16935_/Q vssd1 vssd1 vccd1 vccd1 hold3382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold3393 _11326_/X vssd1 vssd1 vccd1 vccd1 _16932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__buf_4
Xhold2670 _17781_/Q vssd1 vssd1 vccd1 vccd1 hold2670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ hold1746/X _14882_/B _14850_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14851_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2681 _15651_/Q vssd1 vssd1 vccd1 vccd1 hold2681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2692 _14579_/X vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _17721_/Q _13805_/B _13805_/C vssd1 vssd1 vccd1 vccd1 _13802_/X sky130_fd_sc_hd__and3_1
X_17570_ _17730_/CLK _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1980 _14223_/X vssd1 vssd1 vccd1 vccd1 _17913_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14782_ _15229_/A _14786_/B vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__or2_1
Xhold1991 _08226_/X vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ _12282_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__or2_1
X_16521_ _18319_/CLK _16521_/D vssd1 vssd1 vccd1 vccd1 _16521_/Q sky130_fd_sc_hd__dfxtp_1
X_13733_ hold1634/X hold4283/X _13829_/C vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__mux2_1
X_10945_ hold5411/X _11156_/B _10944_/X _14907_/C1 vssd1 vssd1 vccd1 vccd1 _10945_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_45_wb_clk_i clkbuf_leaf_47_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18461_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16452_ _18399_/CLK _16452_/D vssd1 vssd1 vccd1 vccd1 _16452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ hold2842/X hold4641/X _13865_/C vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10876_ hold3948/X _11201_/B _10875_/X _15036_/A vssd1 vssd1 vccd1 vccd1 _10876_/X
+ sky130_fd_sc_hd__o211a_1
X_15403_ _15481_/A1 _15395_/X _15402_/X _15481_/B1 _18416_/Q vssd1 vssd1 vccd1 vccd1
+ _15403_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12924_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _17381_/D sky130_fd_sc_hd__and2_1
X_16383_ _18392_/CLK _16383_/D vssd1 vssd1 vccd1 vccd1 _16383_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13595_ hold2830/X hold5203/X _13883_/C vssd1 vssd1 vccd1 vccd1 _13596_/B sky130_fd_sc_hd__mux2_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _18218_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_1
X_15334_ _15334_/A _15334_/B vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__and2_1
X_12546_ _12933_/A _12546_/B vssd1 vssd1 vccd1 vccd1 _17358_/D sky130_fd_sc_hd__and2_1
XFILLER_0_164_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18053_ _18053_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15265_ hold579/X _15483_/B vssd1 vssd1 vccd1 vccd1 _15265_/X sky130_fd_sc_hd__or2_1
X_12477_ hold11/X _08598_/B _08999_/B _12476_/X _15284_/A vssd1 vssd1 vccd1 vccd1
+ hold12/A sky130_fd_sc_hd__o311a_1
XFILLER_0_112_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17004_ _17852_/CLK _17004_/D vssd1 vssd1 vccd1 vccd1 _17004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_4 _13308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14897_/A hold273/X vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nor2_2
X_11428_ hold5070/X _12305_/B _11427_/X _14149_/C1 vssd1 vssd1 vccd1 vccd1 _11428_/X
+ sky130_fd_sc_hd__o211a_1
X_15196_ hold5967/X _15219_/B hold1342/X _15050_/A vssd1 vssd1 vccd1 vccd1 _15196_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14147_ hold2042/X _14148_/B _14146_/Y _14147_/C1 vssd1 vssd1 vccd1 vccd1 _14147_/X
+ sky130_fd_sc_hd__o211a_1
X_11359_ hold3408/X _12323_/B _11358_/X _13909_/A vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o211a_1
X_14078_ _15531_/A _14106_/B vssd1 vssd1 vccd1 vccd1 _14078_/X sky130_fd_sc_hd__or2_1
X_13029_ _13030_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _17906_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_1
X_17837_ _17892_/CLK hold992/X vssd1 vssd1 vccd1 vccd1 hold991/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ hold17/X hold89/X _08590_/S vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17768_ _17903_/CLK _17768_/D vssd1 vssd1 vccd1 vccd1 _17768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _18020_/CLK _16719_/D vssd1 vssd1 vccd1 vccd1 _16719_/Q sky130_fd_sc_hd__dfxtp_1
X_17699_ _17731_/CLK _17699_/D vssd1 vssd1 vccd1 vccd1 _17699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09122_ _09122_/A hold801/X vssd1 vssd1 vccd1 vccd1 hold802/A sky130_fd_sc_hd__nor2_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09053_ _15354_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _16143_/D sky130_fd_sc_hd__and2_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08004_ hold1136/X _08033_/B _08003_/X _08153_/A vssd1 vssd1 vccd1 vccd1 _08004_/X
+ sky130_fd_sc_hd__o211a_1
Xhold510 hold510/A vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold532 hold532/A vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 hold543/A vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 hold554/A vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold576/A vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 hold587/A vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__clkbuf_8
Xhold598 hold598/A vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ hold5160/X _10049_/B _09954_/X _15070_/A vssd1 vssd1 vccd1 vccd1 _09955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08906_ hold219/X hold696/X _08930_/S vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__mux2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ hold4484/X _10022_/B _09885_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _09886_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _15858_/Q vssd1 vssd1 vccd1 vccd1 hold1210/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _14933_/X vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1232 _07955_/X vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _13002_/A _08837_/B vssd1 vssd1 vccd1 vccd1 _16037_/D sky130_fd_sc_hd__and2_1
Xhold1243 _08286_/X vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1254 _14073_/X vssd1 vssd1 vccd1 vccd1 _17841_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1265 _17844_/Q vssd1 vssd1 vccd1 vccd1 hold1265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 _08294_/X vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _15146_/X vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _15354_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _16004_/D sky130_fd_sc_hd__and2_1
Xhold1298 input59/X vssd1 vssd1 vccd1 vccd1 hold1298/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ hold184/X hold702/X _08721_/S vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ hold2285/X hold3601/X _11762_/C vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ _17914_/Q hold3610/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_137_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12400_ _13002_/A _12400_/B vssd1 vssd1 vccd1 vccd1 _17293_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ _13764_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__or2_1
X_10592_ _10592_/A _10646_/B _10646_/C vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__and3_1
XFILLER_0_134_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _12331_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_163_wb_clk_i clkbuf_5_31__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18192_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15050_ _15050_/A _15050_/B vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12262_ hold4961/X _12356_/B _12261_/X _08139_/A vssd1 vssd1 vccd1 vccd1 _12262_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _14681_/A hold272/X vssd1 vssd1 vccd1 vccd1 _14050_/B sky130_fd_sc_hd__or2_4
X_11213_ _16895_/Q _11213_/B _11213_/C vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__and3_1
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ hold4217/X _12308_/B _12192_/X _08163_/A vssd1 vssd1 vccd1 vccd1 _17221_/D
+ sky130_fd_sc_hd__o211a_1
X_11144_ _16872_/Q _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11144_/X sky130_fd_sc_hd__and3_1
Xoutput74 _13145_/A vssd1 vssd1 vccd1 vccd1 output74/X sky130_fd_sc_hd__buf_6
Xoutput85 _13225_/A vssd1 vssd1 vccd1 vccd1 output85/X sky130_fd_sc_hd__buf_6
Xoutput96 _13305_/A vssd1 vssd1 vccd1 vccd1 output96/X sky130_fd_sc_hd__buf_6
XFILLER_0_179_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15952_ _17342_/CLK _15952_/D vssd1 vssd1 vccd1 vccd1 hold531/A sky130_fd_sc_hd__dfxtp_1
X_11075_ hold971/X hold3299/X _11171_/C vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3190 _10570_/Y vssd1 vssd1 vccd1 vccd1 _16680_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10026_ _13182_/A _09924_/A _10025_/X vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__a21oi_1
X_14903_ hold1927/X hold657/A _14902_/X _15032_/A vssd1 vssd1 vccd1 vccd1 _14903_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15883_ _17723_/CLK _15883_/D vssd1 vssd1 vccd1 vccd1 _15883_/Q sky130_fd_sc_hd__dfxtp_1
X_17622_ _17686_/CLK _17622_/D vssd1 vssd1 vccd1 vccd1 _17622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14834_ _15227_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _18229_/CLK _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ hold2730/X _14774_/B _14764_/X _14863_/C1 vssd1 vssd1 vccd1 vccd1 _14765_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ hold5112/X _13871_/B _11976_/X _08141_/A vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _18385_/CLK _16504_/D vssd1 vssd1 vccd1 vccd1 _16504_/Q sky130_fd_sc_hd__dfxtp_1
X_13716_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__or2_1
X_17484_ _17484_/CLK _17484_/D vssd1 vssd1 vccd1 vccd1 _17484_/Q sky130_fd_sc_hd__dfxtp_1
X_10928_ hold1294/X hold5518/X _11216_/C vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__mux2_1
X_14696_ _15197_/A _14732_/B vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16435_ _18386_/CLK _16435_/D vssd1 vssd1 vccd1 vccd1 _16435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13776_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__or2_1
X_10859_ hold2456/X hold3240/X _11153_/C vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16366_ _18424_/CLK _16366_/D vssd1 vssd1 vccd1 vccd1 _16366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13674_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__or2_1
X_18105_ _18149_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15317_ hold287/X _09357_/A _15484_/B1 hold338/X _15316_/X vssd1 vssd1 vccd1 vccd1
+ _15322_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ hold1883/X hold3438/X _13000_/S vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__mux2_1
X_16297_ _17511_/CLK _16297_/D vssd1 vssd1 vccd1 vccd1 _16297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5509 _10861_/X vssd1 vssd1 vccd1 vccd1 _16777_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _18070_/CLK hold790/X vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ hold409/X _15484_/A2 _15451_/A2 hold473/X vssd1 vssd1 vccd1 vccd1 _15248_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4808 _13711_/X vssd1 vssd1 vccd1 vccd1 _17690_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4819 _11959_/X vssd1 vssd1 vccd1 vccd1 _17143_/D sky130_fd_sc_hd__dlygate4sd3_1
X_15179_ _15233_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__or2_1
Xfanout308 _09918_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__buf_4
Xfanout319 _10998_/A vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__buf_4
X_09740_ hold1477/X _16404_/Q _10067_/C vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

