VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vmsu_8bit_top
  CLASS BLOCK ;
  FOREIGN vmsu_8bit_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END b[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clk
  PIN control
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END control
  PIN p[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END p[15]
  PIN p[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 485.465 494.230 487.070 ;
        RECT 5.330 480.025 494.230 482.855 ;
        RECT 5.330 474.585 494.230 477.415 ;
        RECT 5.330 469.145 494.230 471.975 ;
        RECT 5.330 463.705 494.230 466.535 ;
        RECT 5.330 458.265 494.230 461.095 ;
        RECT 5.330 452.825 494.230 455.655 ;
        RECT 5.330 447.385 494.230 450.215 ;
        RECT 5.330 441.945 494.230 444.775 ;
        RECT 5.330 436.505 494.230 439.335 ;
        RECT 5.330 431.065 494.230 433.895 ;
        RECT 5.330 425.625 494.230 428.455 ;
        RECT 5.330 420.185 494.230 423.015 ;
        RECT 5.330 414.745 494.230 417.575 ;
        RECT 5.330 409.305 494.230 412.135 ;
        RECT 5.330 403.865 494.230 406.695 ;
        RECT 5.330 398.425 494.230 401.255 ;
        RECT 5.330 392.985 494.230 395.815 ;
        RECT 5.330 387.545 494.230 390.375 ;
        RECT 5.330 382.105 494.230 384.935 ;
        RECT 5.330 376.665 494.230 379.495 ;
        RECT 5.330 371.225 494.230 374.055 ;
        RECT 5.330 365.785 494.230 368.615 ;
        RECT 5.330 360.345 494.230 363.175 ;
        RECT 5.330 354.905 494.230 357.735 ;
        RECT 5.330 349.465 494.230 352.295 ;
        RECT 5.330 344.025 494.230 346.855 ;
        RECT 5.330 338.585 494.230 341.415 ;
        RECT 5.330 333.145 494.230 335.975 ;
        RECT 5.330 327.705 494.230 330.535 ;
        RECT 5.330 322.265 494.230 325.095 ;
        RECT 5.330 316.825 494.230 319.655 ;
        RECT 5.330 311.385 494.230 314.215 ;
        RECT 5.330 305.945 494.230 308.775 ;
        RECT 5.330 300.505 494.230 303.335 ;
        RECT 5.330 295.065 494.230 297.895 ;
        RECT 5.330 289.625 494.230 292.455 ;
        RECT 5.330 284.185 494.230 287.015 ;
        RECT 5.330 278.745 494.230 281.575 ;
        RECT 5.330 273.305 494.230 276.135 ;
        RECT 5.330 267.865 494.230 270.695 ;
        RECT 5.330 262.425 494.230 265.255 ;
        RECT 5.330 256.985 494.230 259.815 ;
        RECT 5.330 251.545 494.230 254.375 ;
        RECT 5.330 246.105 494.230 248.935 ;
        RECT 5.330 240.665 494.230 243.495 ;
        RECT 5.330 235.225 494.230 238.055 ;
        RECT 5.330 229.785 494.230 232.615 ;
        RECT 5.330 224.345 494.230 227.175 ;
        RECT 5.330 218.905 494.230 221.735 ;
        RECT 5.330 213.465 494.230 216.295 ;
        RECT 5.330 208.025 494.230 210.855 ;
        RECT 5.330 202.585 494.230 205.415 ;
        RECT 5.330 197.145 494.230 199.975 ;
        RECT 5.330 191.705 494.230 194.535 ;
        RECT 5.330 186.265 494.230 189.095 ;
        RECT 5.330 180.825 494.230 183.655 ;
        RECT 5.330 175.385 494.230 178.215 ;
        RECT 5.330 169.945 494.230 172.775 ;
        RECT 5.330 164.505 494.230 167.335 ;
        RECT 5.330 159.065 494.230 161.895 ;
        RECT 5.330 153.625 494.230 156.455 ;
        RECT 5.330 148.185 494.230 151.015 ;
        RECT 5.330 142.745 494.230 145.575 ;
        RECT 5.330 137.305 494.230 140.135 ;
        RECT 5.330 131.865 494.230 134.695 ;
        RECT 5.330 126.425 494.230 129.255 ;
        RECT 5.330 120.985 494.230 123.815 ;
        RECT 5.330 115.545 494.230 118.375 ;
        RECT 5.330 110.105 494.230 112.935 ;
        RECT 5.330 104.665 494.230 107.495 ;
        RECT 5.330 99.225 494.230 102.055 ;
        RECT 5.330 93.785 494.230 96.615 ;
        RECT 5.330 88.345 494.230 91.175 ;
        RECT 5.330 82.905 494.230 85.735 ;
        RECT 5.330 77.465 494.230 80.295 ;
        RECT 5.330 72.025 494.230 74.855 ;
        RECT 5.330 66.585 494.230 69.415 ;
        RECT 5.330 61.145 494.230 63.975 ;
        RECT 5.330 55.705 494.230 58.535 ;
        RECT 5.330 50.265 494.230 53.095 ;
        RECT 5.330 44.825 494.230 47.655 ;
        RECT 5.330 39.385 494.230 42.215 ;
        RECT 5.330 33.945 494.230 36.775 ;
        RECT 5.330 28.505 494.230 31.335 ;
        RECT 5.330 23.065 494.230 25.895 ;
        RECT 5.330 17.625 494.230 20.455 ;
        RECT 5.330 12.185 494.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 7.460 4.280 492.500 487.065 ;
        RECT 8.010 3.670 21.430 4.280 ;
        RECT 22.270 3.670 35.690 4.280 ;
        RECT 36.530 3.670 49.950 4.280 ;
        RECT 50.790 3.670 64.210 4.280 ;
        RECT 65.050 3.670 78.470 4.280 ;
        RECT 79.310 3.670 92.730 4.280 ;
        RECT 93.570 3.670 106.990 4.280 ;
        RECT 107.830 3.670 121.250 4.280 ;
        RECT 122.090 3.670 135.510 4.280 ;
        RECT 136.350 3.670 149.770 4.280 ;
        RECT 150.610 3.670 164.030 4.280 ;
        RECT 164.870 3.670 178.290 4.280 ;
        RECT 179.130 3.670 192.550 4.280 ;
        RECT 193.390 3.670 206.810 4.280 ;
        RECT 207.650 3.670 221.070 4.280 ;
        RECT 221.910 3.670 235.330 4.280 ;
        RECT 236.170 3.670 249.590 4.280 ;
        RECT 250.430 3.670 263.850 4.280 ;
        RECT 264.690 3.670 278.110 4.280 ;
        RECT 278.950 3.670 292.370 4.280 ;
        RECT 293.210 3.670 306.630 4.280 ;
        RECT 307.470 3.670 320.890 4.280 ;
        RECT 321.730 3.670 335.150 4.280 ;
        RECT 335.990 3.670 349.410 4.280 ;
        RECT 350.250 3.670 363.670 4.280 ;
        RECT 364.510 3.670 377.930 4.280 ;
        RECT 378.770 3.670 392.190 4.280 ;
        RECT 393.030 3.670 406.450 4.280 ;
        RECT 407.290 3.670 420.710 4.280 ;
        RECT 421.550 3.670 434.970 4.280 ;
        RECT 435.810 3.670 449.230 4.280 ;
        RECT 450.070 3.670 463.490 4.280 ;
        RECT 464.330 3.670 477.750 4.280 ;
        RECT 478.590 3.670 492.010 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 483.430 487.045 ;
  END
END vmsu_8bit_top
END LIBRARY

